`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper : Time Sharing - A Novel Approach to Low-Latency Masking
// Authors : Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date:    00:33:45 09/30/2023 
// Design Name:    AES S-Box 
// Module Name:    AES_sbox_opt 
// Description:    Top module for AES S-Box.  
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module AES_sbox_opt (clk, PRNG_rand, sbox_input_share1, sbox_input_share2,  sbox_output_share1, sbox_output_share2);

input clk ;
input [262:1] PRNG_rand ; 
input [7:0] sbox_input_share1, sbox_input_share2 ;
output [7:0] sbox_output_share1, sbox_output_share2 ;

wire [7:0] rand_composable_bit ;

assign rand_composable_bit = PRNG_rand[8:1] ;

reg x0_subscript0_share1_reg , x2_subscript0_share1_reg , x3_subscript0_share1_reg , x4_subscript0_share1_reg , x6_subscript0_share1_reg , x7_subscript0_share1_reg , x1_subscript0_share1_reg , x5_subscript0_share1_reg , x0x1_subscript0_share1_reg , x0x4_subscript0_share1_reg , x0x5_subscript0_share1_reg , x0x6_subscript0_share1_reg , x1x2_subscript0_share1_reg , x1x3_subscript0_share1_reg , x1x4_subscript0_share1_reg , x1x6_subscript0_share1_reg , x2x3_subscript0_share1_reg , x2x4_subscript0_share1_reg , x2x6_subscript0_share1_reg , x2x7_subscript0_share1_reg , x4x6_subscript0_share1_reg , x5x6_subscript0_share1_reg , x5x7_subscript0_share1_reg , x6x7_subscript0_share1_reg , x0x2_subscript0_share1_reg , x0x3_subscript0_share1_reg , x0x7_subscript0_share1_reg , x1x7_subscript0_share1_reg , x3x7_subscript0_share1_reg , x4x5_subscript0_share1_reg , x3x4_subscript0_share1_reg , x4x7_subscript0_share1_reg , x3x6_subscript0_share1_reg , x1x5_subscript0_share1_reg , x2x5_subscript0_share1_reg , x3x5_subscript0_share1_reg , x0x1x4_subscript0_share1_reg , x0x1x6_subscript0_share1_reg , x0x1x7_subscript0_share1_reg , x0x2x4_subscript0_share1_reg , x0x2x5_subscript0_share1_reg , x0x2x6_subscript0_share1_reg , x0x2x7_subscript0_share1_reg , x0x3x4_subscript0_share1_reg , x0x3x5_subscript0_share1_reg , x0x3x6_subscript0_share1_reg , x0x4x6_subscript0_share1_reg , x0x4x7_subscript0_share1_reg , x1x2x3_subscript0_share1_reg , x1x2x4_subscript0_share1_reg , x1x2x6_subscript0_share1_reg , x1x3x4_subscript0_share1_reg , x1x3x7_subscript0_share1_reg , x1x4x6_subscript0_share1_reg , x1x5x6_subscript0_share1_reg , x2x3x5_subscript0_share1_reg , x2x3x7_subscript0_share1_reg , x2x4x7_subscript0_share1_reg , x2x5x6_subscript0_share1_reg , x2x5x7_subscript0_share1_reg , x2x6x7_subscript0_share1_reg , x3x4x7_subscript0_share1_reg , x3x5x7_subscript0_share1_reg , x3x6x7_subscript0_share1_reg , x4x5x6_subscript0_share1_reg , x5x6x7_subscript0_share1_reg , x0x1x3_subscript0_share1_reg , x0x2x3_subscript0_share1_reg , x0x4x5_subscript0_share1_reg , x0x5x7_subscript0_share1_reg , x0x6x7_subscript0_share1_reg , x1x3x5_subscript0_share1_reg , x1x3x6_subscript0_share1_reg , x1x4x7_subscript0_share1_reg , x2x3x4_subscript0_share1_reg , x2x3x6_subscript0_share1_reg , x3x4x6_subscript0_share1_reg , x3x5x6_subscript0_share1_reg , x0x1x5_subscript0_share1_reg , x0x3x7_subscript0_share1_reg , x1x2x5_subscript0_share1_reg , x1x2x7_subscript0_share1_reg , x1x4x5_subscript0_share1_reg , x1x5x7_subscript0_share1_reg , x2x4x5_subscript0_share1_reg , x3x4x5_subscript0_share1_reg , x4x6x7_subscript0_share1_reg , x1x6x7_subscript0_share1_reg , x4x5x7_subscript0_share1_reg , x0x1x2_subscript0_share1_reg , x0x5x6_subscript0_share1_reg , x2x4x6_subscript0_share1_reg , x0x1x2x3_subscript0_share1_reg , x0x1x2x5_subscript0_share1_reg , x0x1x2x6_subscript0_share1_reg , x0x1x2x7_subscript0_share1_reg , x0x1x4x5_subscript0_share1_reg , x0x1x4x7_subscript0_share1_reg , x0x2x3x5_subscript0_share1_reg , x0x2x3x7_subscript0_share1_reg , x0x2x4x5_subscript0_share1_reg , x0x2x4x7_subscript0_share1_reg , x0x2x5x6_subscript0_share1_reg , x0x2x5x7_subscript0_share1_reg , x0x3x4x6_subscript0_share1_reg , x0x3x5x6_subscript0_share1_reg , x0x4x5x6_subscript0_share1_reg , x0x4x5x7_subscript0_share1_reg , x0x4x6x7_subscript0_share1_reg , x1x2x3x5_subscript0_share1_reg , x1x2x3x6_subscript0_share1_reg , x1x2x3x7_subscript0_share1_reg , x1x2x4x6_subscript0_share1_reg , x1x2x4x7_subscript0_share1_reg , x1x2x6x7_subscript0_share1_reg , x1x3x4x6_subscript0_share1_reg , x1x3x6x7_subscript0_share1_reg , x1x4x5x6_subscript0_share1_reg , x1x4x5x7_subscript0_share1_reg , x1x5x6x7_subscript0_share1_reg , x2x3x5x7_subscript0_share1_reg , x2x3x6x7_subscript0_share1_reg , x2x4x5x6_subscript0_share1_reg , x2x4x5x7_subscript0_share1_reg , x3x5x6x7_subscript0_share1_reg , x0x1x3x4_subscript0_share1_reg , x0x1x3x6_subscript0_share1_reg , x0x1x5x6_subscript0_share1_reg , x0x2x3x6_subscript0_share1_reg , x0x3x4x5_subscript0_share1_reg , x1x2x5x6_subscript0_share1_reg , x1x2x5x7_subscript0_share1_reg , x1x3x4x5_subscript0_share1_reg , x1x3x4x7_subscript0_share1_reg , x1x3x5x6_subscript0_share1_reg , x1x3x5x7_subscript0_share1_reg , x1x4x6x7_subscript0_share1_reg , x2x3x4x5_subscript0_share1_reg , x2x3x4x7_subscript0_share1_reg , x2x4x6x7_subscript0_share1_reg , x3x4x5x6_subscript0_share1_reg , x3x4x5x7_subscript0_share1_reg , x3x4x6x7_subscript0_share1_reg , x0x1x3x5_subscript0_share1_reg , x0x1x4x6_subscript0_share1_reg , x0x2x3x4_subscript0_share1_reg , x0x2x4x6_subscript0_share1_reg , x0x3x4x7_subscript0_share1_reg , x0x3x5x7_subscript0_share1_reg , x1x2x3x4_subscript0_share1_reg , x2x3x4x6_subscript0_share1_reg , x2x3x5x6_subscript0_share1_reg , x2x5x6x7_subscript0_share1_reg , x4x5x6x7_subscript0_share1_reg , x0x1x2x4_subscript0_share1_reg , x0x1x6x7_subscript0_share1_reg , x0x2x6x7_subscript0_share1_reg , x0x3x6x7_subscript0_share1_reg , x0x5x6x7_subscript0_share1_reg , x1x2x4x5_subscript0_share1_reg , x0x1x3x7_subscript0_share1_reg , x0x1x5x7_subscript0_share1_reg , x0x1x2x3x4_subscript0_share1_reg , x0x1x2x3x6_subscript0_share1_reg , x0x1x2x3x7_subscript0_share1_reg , x0x1x2x4x5_subscript0_share1_reg , x0x1x2x4x7_subscript0_share1_reg , x0x1x2x5x7_subscript0_share1_reg , x0x1x2x6x7_subscript0_share1_reg , x0x1x3x4x6_subscript0_share1_reg , x0x1x3x5x6_subscript0_share1_reg , x0x1x3x5x7_subscript0_share1_reg , x0x1x3x6x7_subscript0_share1_reg , x0x1x4x5x6_subscript0_share1_reg , x0x1x5x6x7_subscript0_share1_reg , x0x2x3x4x5_subscript0_share1_reg , x0x2x3x4x6_subscript0_share1_reg , x0x2x4x5x7_subscript0_share1_reg , x0x2x4x6x7_subscript0_share1_reg , x0x3x4x5x6_subscript0_share1_reg , x0x3x4x5x7_subscript0_share1_reg , x0x3x4x6x7_subscript0_share1_reg , x0x3x5x6x7_subscript0_share1_reg , x1x2x3x5x6_subscript0_share1_reg , x1x2x3x5x7_subscript0_share1_reg , x1x2x4x5x6_subscript0_share1_reg , x1x2x4x6x7_subscript0_share1_reg , x1x2x5x6x7_subscript0_share1_reg , x1x3x4x5x7_subscript0_share1_reg , x2x3x4x5x6_subscript0_share1_reg , x2x3x4x5x7_subscript0_share1_reg , x2x4x5x6x7_subscript0_share1_reg , x0x1x2x4x6_subscript0_share1_reg , x0x1x3x4x7_subscript0_share1_reg , x0x2x3x4x7_subscript0_share1_reg , x0x2x3x5x7_subscript0_share1_reg , x0x2x3x6x7_subscript0_share1_reg , x0x2x4x5x6_subscript0_share1_reg , x0x2x5x6x7_subscript0_share1_reg , x0x4x5x6x7_subscript0_share1_reg , x1x2x3x4x6_subscript0_share1_reg , x1x3x4x5x6_subscript0_share1_reg , x2x3x4x6x7_subscript0_share1_reg , x0x1x2x3x5_subscript0_share1_reg , x0x1x4x6x7_subscript0_share1_reg , x1x2x3x4x5_subscript0_share1_reg , x1x2x3x6x7_subscript0_share1_reg , x1x2x4x5x7_subscript0_share1_reg , x1x3x4x6x7_subscript0_share1_reg , x1x3x5x6x7_subscript0_share1_reg , x1x4x5x6x7_subscript0_share1_reg , x2x3x5x6x7_subscript0_share1_reg , x3x4x5x6x7_subscript0_share1_reg , x0x1x2x5x6_subscript0_share1_reg , x0x1x3x4x5_subscript0_share1_reg , x0x1x4x5x7_subscript0_share1_reg , x0x2x3x5x6_subscript0_share1_reg , x1x2x3x4x7_subscript0_share1_reg , x0x1x2x3x4x6_subscript0_share1_reg , x0x1x2x3x4x7_subscript0_share1_reg , x0x1x2x3x5x7_subscript0_share1_reg , x0x1x2x3x6x7_subscript0_share1_reg , x0x1x2x4x5x7_subscript0_share1_reg , x0x1x2x5x6x7_subscript0_share1_reg , x0x1x3x4x6x7_subscript0_share1_reg , x0x1x4x5x6x7_subscript0_share1_reg , x0x2x3x4x5x6_subscript0_share1_reg , x0x2x3x4x5x7_subscript0_share1_reg , x0x2x3x5x6x7_subscript0_share1_reg , x1x2x3x4x6x7_subscript0_share1_reg , x1x2x4x5x6x7_subscript0_share1_reg , x1x3x4x5x6x7_subscript0_share1_reg , x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x5x6_subscript0_share1_reg , x0x1x2x4x6x7_subscript0_share1_reg , x0x1x3x4x5x6_subscript0_share1_reg , x0x2x3x4x6x7_subscript0_share1_reg , x1x2x3x4x5x6_subscript0_share1_reg , x1x2x3x5x6x7_subscript0_share1_reg , x0x1x2x3x4x5_subscript0_share1_reg , x0x1x2x4x5x6_subscript0_share1_reg , x0x1x3x4x5x7_subscript0_share1_reg , x0x1x3x5x6x7_subscript0_share1_reg , x0x2x4x5x6x7_subscript0_share1_reg , x1x2x3x4x5x7_subscript0_share1_reg , x0x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x4x6x7_subscript0_share1_reg , x0x1x2x4x5x6x7_subscript0_share1_reg , x0x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x5x6x7_subscript0_share1_reg , x0x1x3x4x5x6x7_subscript0_share1_reg , x1x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x4x5x6_subscript0_share1_reg , x0x1x2x3x4x5x7_subscript0_share1_reg ;
reg x0_subscript0_share2_reg , x2_subscript0_share2_reg , x3_subscript0_share2_reg , x4_subscript0_share2_reg , x6_subscript0_share2_reg , x7_subscript0_share2_reg , x1_subscript0_share2_reg , x5_subscript0_share2_reg , x0x1_subscript0_share2_reg , x0x4_subscript0_share2_reg , x0x5_subscript0_share2_reg , x0x6_subscript0_share2_reg , x1x2_subscript0_share2_reg , x1x3_subscript0_share2_reg , x1x4_subscript0_share2_reg , x1x6_subscript0_share2_reg , x2x3_subscript0_share2_reg , x2x4_subscript0_share2_reg , x2x6_subscript0_share2_reg , x2x7_subscript0_share2_reg , x4x6_subscript0_share2_reg , x5x6_subscript0_share2_reg , x5x7_subscript0_share2_reg , x6x7_subscript0_share2_reg , x0x2_subscript0_share2_reg , x0x3_subscript0_share2_reg , x0x7_subscript0_share2_reg , x1x7_subscript0_share2_reg , x3x7_subscript0_share2_reg , x4x5_subscript0_share2_reg , x3x4_subscript0_share2_reg , x4x7_subscript0_share2_reg , x3x6_subscript0_share2_reg , x1x5_subscript0_share2_reg , x2x5_subscript0_share2_reg , x3x5_subscript0_share2_reg , x0x1x4_subscript0_share2_reg , x0x1x6_subscript0_share2_reg , x0x1x7_subscript0_share2_reg , x0x2x4_subscript0_share2_reg , x0x2x5_subscript0_share2_reg , x0x2x6_subscript0_share2_reg , x0x2x7_subscript0_share2_reg , x0x3x4_subscript0_share2_reg , x0x3x5_subscript0_share2_reg , x0x3x6_subscript0_share2_reg , x0x4x6_subscript0_share2_reg , x0x4x7_subscript0_share2_reg , x1x2x3_subscript0_share2_reg , x1x2x4_subscript0_share2_reg , x1x2x6_subscript0_share2_reg , x1x3x4_subscript0_share2_reg , x1x3x7_subscript0_share2_reg , x1x4x6_subscript0_share2_reg , x1x5x6_subscript0_share2_reg , x2x3x5_subscript0_share2_reg , x2x3x7_subscript0_share2_reg , x2x4x7_subscript0_share2_reg , x2x5x6_subscript0_share2_reg , x2x5x7_subscript0_share2_reg , x2x6x7_subscript0_share2_reg , x3x4x7_subscript0_share2_reg , x3x5x7_subscript0_share2_reg , x3x6x7_subscript0_share2_reg , x4x5x6_subscript0_share2_reg , x5x6x7_subscript0_share2_reg , x0x1x3_subscript0_share2_reg , x0x2x3_subscript0_share2_reg , x0x4x5_subscript0_share2_reg , x0x5x7_subscript0_share2_reg , x0x6x7_subscript0_share2_reg , x1x3x5_subscript0_share2_reg , x1x3x6_subscript0_share2_reg , x1x4x7_subscript0_share2_reg , x2x3x4_subscript0_share2_reg , x2x3x6_subscript0_share2_reg , x3x4x6_subscript0_share2_reg , x3x5x6_subscript0_share2_reg , x0x1x5_subscript0_share2_reg , x0x3x7_subscript0_share2_reg , x1x2x5_subscript0_share2_reg , x1x2x7_subscript0_share2_reg , x1x4x5_subscript0_share2_reg , x1x5x7_subscript0_share2_reg , x2x4x5_subscript0_share2_reg , x3x4x5_subscript0_share2_reg , x4x6x7_subscript0_share2_reg , x1x6x7_subscript0_share2_reg , x4x5x7_subscript0_share2_reg , x0x1x2_subscript0_share2_reg , x0x5x6_subscript0_share2_reg , x2x4x6_subscript0_share2_reg , x0x1x2x3_subscript0_share2_reg , x0x1x2x5_subscript0_share2_reg , x0x1x2x6_subscript0_share2_reg , x0x1x2x7_subscript0_share2_reg , x0x1x4x5_subscript0_share2_reg , x0x1x4x7_subscript0_share2_reg , x0x2x3x5_subscript0_share2_reg , x0x2x3x7_subscript0_share2_reg , x0x2x4x5_subscript0_share2_reg , x0x2x4x7_subscript0_share2_reg , x0x2x5x6_subscript0_share2_reg , x0x2x5x7_subscript0_share2_reg , x0x3x4x6_subscript0_share2_reg , x0x3x5x6_subscript0_share2_reg , x0x4x5x6_subscript0_share2_reg , x0x4x5x7_subscript0_share2_reg , x0x4x6x7_subscript0_share2_reg , x1x2x3x5_subscript0_share2_reg , x1x2x3x6_subscript0_share2_reg , x1x2x3x7_subscript0_share2_reg , x1x2x4x6_subscript0_share2_reg , x1x2x4x7_subscript0_share2_reg , x1x2x6x7_subscript0_share2_reg , x1x3x4x6_subscript0_share2_reg , x1x3x6x7_subscript0_share2_reg , x1x4x5x6_subscript0_share2_reg , x1x4x5x7_subscript0_share2_reg , x1x5x6x7_subscript0_share2_reg , x2x3x5x7_subscript0_share2_reg , x2x3x6x7_subscript0_share2_reg , x2x4x5x6_subscript0_share2_reg , x2x4x5x7_subscript0_share2_reg , x3x5x6x7_subscript0_share2_reg , x0x1x3x4_subscript0_share2_reg , x0x1x3x6_subscript0_share2_reg , x0x1x5x6_subscript0_share2_reg , x0x2x3x6_subscript0_share2_reg , x0x3x4x5_subscript0_share2_reg , x1x2x5x6_subscript0_share2_reg , x1x2x5x7_subscript0_share2_reg , x1x3x4x5_subscript0_share2_reg , x1x3x4x7_subscript0_share2_reg , x1x3x5x6_subscript0_share2_reg , x1x3x5x7_subscript0_share2_reg , x1x4x6x7_subscript0_share2_reg , x2x3x4x5_subscript0_share2_reg , x2x3x4x7_subscript0_share2_reg , x2x4x6x7_subscript0_share2_reg , x3x4x5x6_subscript0_share2_reg , x3x4x5x7_subscript0_share2_reg , x3x4x6x7_subscript0_share2_reg , x0x1x3x5_subscript0_share2_reg , x0x1x4x6_subscript0_share2_reg , x0x2x3x4_subscript0_share2_reg , x0x2x4x6_subscript0_share2_reg , x0x3x4x7_subscript0_share2_reg , x0x3x5x7_subscript0_share2_reg , x1x2x3x4_subscript0_share2_reg , x2x3x4x6_subscript0_share2_reg , x2x3x5x6_subscript0_share2_reg , x2x5x6x7_subscript0_share2_reg , x4x5x6x7_subscript0_share2_reg , x0x1x2x4_subscript0_share2_reg , x0x1x6x7_subscript0_share2_reg , x0x2x6x7_subscript0_share2_reg , x0x3x6x7_subscript0_share2_reg , x0x5x6x7_subscript0_share2_reg , x1x2x4x5_subscript0_share2_reg , x0x1x3x7_subscript0_share2_reg , x0x1x5x7_subscript0_share2_reg , x0x1x2x3x4_subscript0_share2_reg , x0x1x2x3x6_subscript0_share2_reg , x0x1x2x3x7_subscript0_share2_reg , x0x1x2x4x5_subscript0_share2_reg , x0x1x2x4x7_subscript0_share2_reg , x0x1x2x5x7_subscript0_share2_reg , x0x1x2x6x7_subscript0_share2_reg , x0x1x3x4x6_subscript0_share2_reg , x0x1x3x5x6_subscript0_share2_reg , x0x1x3x5x7_subscript0_share2_reg , x0x1x3x6x7_subscript0_share2_reg , x0x1x4x5x6_subscript0_share2_reg , x0x1x5x6x7_subscript0_share2_reg , x0x2x3x4x5_subscript0_share2_reg , x0x2x3x4x6_subscript0_share2_reg , x0x2x4x5x7_subscript0_share2_reg , x0x2x4x6x7_subscript0_share2_reg , x0x3x4x5x6_subscript0_share2_reg , x0x3x4x5x7_subscript0_share2_reg , x0x3x4x6x7_subscript0_share2_reg , x0x3x5x6x7_subscript0_share2_reg , x1x2x3x5x6_subscript0_share2_reg , x1x2x3x5x7_subscript0_share2_reg , x1x2x4x5x6_subscript0_share2_reg , x1x2x4x6x7_subscript0_share2_reg , x1x2x5x6x7_subscript0_share2_reg , x1x3x4x5x7_subscript0_share2_reg , x2x3x4x5x6_subscript0_share2_reg , x2x3x4x5x7_subscript0_share2_reg , x2x4x5x6x7_subscript0_share2_reg , x0x1x2x4x6_subscript0_share2_reg , x0x1x3x4x7_subscript0_share2_reg , x0x2x3x4x7_subscript0_share2_reg , x0x2x3x5x7_subscript0_share2_reg , x0x2x3x6x7_subscript0_share2_reg , x0x2x4x5x6_subscript0_share2_reg , x0x2x5x6x7_subscript0_share2_reg , x0x4x5x6x7_subscript0_share2_reg , x1x2x3x4x6_subscript0_share2_reg , x1x3x4x5x6_subscript0_share2_reg , x2x3x4x6x7_subscript0_share2_reg , x0x1x2x3x5_subscript0_share2_reg , x0x1x4x6x7_subscript0_share2_reg , x1x2x3x4x5_subscript0_share2_reg , x1x2x3x6x7_subscript0_share2_reg , x1x2x4x5x7_subscript0_share2_reg , x1x3x4x6x7_subscript0_share2_reg , x1x3x5x6x7_subscript0_share2_reg , x1x4x5x6x7_subscript0_share2_reg , x2x3x5x6x7_subscript0_share2_reg , x3x4x5x6x7_subscript0_share2_reg , x0x1x2x5x6_subscript0_share2_reg , x0x1x3x4x5_subscript0_share2_reg , x0x1x4x5x7_subscript0_share2_reg , x0x2x3x5x6_subscript0_share2_reg , x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x4x6_subscript0_share2_reg , x0x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x5x7_subscript0_share2_reg , x0x1x2x3x6x7_subscript0_share2_reg , x0x1x2x4x5x7_subscript0_share2_reg , x0x1x2x5x6x7_subscript0_share2_reg , x0x1x3x4x6x7_subscript0_share2_reg , x0x1x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6_subscript0_share2_reg , x0x2x3x4x5x7_subscript0_share2_reg , x0x2x3x5x6x7_subscript0_share2_reg , x1x2x3x4x6x7_subscript0_share2_reg , x1x2x4x5x6x7_subscript0_share2_reg , x1x3x4x5x6x7_subscript0_share2_reg , x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6_subscript0_share2_reg , x0x1x2x4x6x7_subscript0_share2_reg , x0x1x3x4x5x6_subscript0_share2_reg , x0x2x3x4x6x7_subscript0_share2_reg , x1x2x3x4x5x6_subscript0_share2_reg , x1x2x3x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5_subscript0_share2_reg , x0x1x2x4x5x6_subscript0_share2_reg , x0x1x3x4x5x7_subscript0_share2_reg , x0x1x3x5x6x7_subscript0_share2_reg , x0x2x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x7_subscript0_share2_reg , x0x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x6x7_subscript0_share2_reg , x0x1x2x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6x7_subscript0_share2_reg , x0x1x3x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5x6_subscript0_share2_reg , x0x1x2x3x4x5x7_subscript0_share2_reg ;
reg x0_share2_reg , x1_share2_reg , x2_share2_reg , x3_share2_reg , x4_share2_reg , x5_share2_reg , x6_share2_reg , x7_share2_reg ;

AES_sbox_compute_subscript0 inst0( sbox_input_share1, PRNG_rand[262:9], rand_composable_bit, x0_subscript0_share1_1 , x2_subscript0_share1_1 , x3_subscript0_share1_1 , x4_subscript0_share1_1 , x6_subscript0_share1_1 , x7_subscript0_share1_1 , x1_subscript0_share1_1 , x5_subscript0_share1_1 , x0x1_subscript0_share1_1 , x0x4_subscript0_share1_1 , x0x5_subscript0_share1_1 , x0x6_subscript0_share1_1 , x1x2_subscript0_share1_1 , x1x3_subscript0_share1_1 , x1x4_subscript0_share1_1 , x1x6_subscript0_share1_1 , x2x3_subscript0_share1_1 , x2x4_subscript0_share1_1 , x2x6_subscript0_share1_1 , x2x7_subscript0_share1_1 , x4x6_subscript0_share1_1 , x5x6_subscript0_share1_1 , x5x7_subscript0_share1_1 , x6x7_subscript0_share1_1 , x0x2_subscript0_share1_1 , x0x3_subscript0_share1_1 , x0x7_subscript0_share1_1 , x1x7_subscript0_share1_1 , x3x7_subscript0_share1_1 , x4x5_subscript0_share1_1 , x3x4_subscript0_share1_1 , x4x7_subscript0_share1_1 , x3x6_subscript0_share1_1 , x1x5_subscript0_share1_1 , x2x5_subscript0_share1_1 , x3x5_subscript0_share1_1 , x0x1x4_subscript0_share1_1 , x0x1x6_subscript0_share1_1 , x0x1x7_subscript0_share1_1 , x0x2x4_subscript0_share1_1 , x0x2x5_subscript0_share1_1 , x0x2x6_subscript0_share1_1 , x0x2x7_subscript0_share1_1 , x0x3x4_subscript0_share1_1 , x0x3x5_subscript0_share1_1 , x0x3x6_subscript0_share1_1 , x0x4x6_subscript0_share1_1 , x0x4x7_subscript0_share1_1 , x1x2x3_subscript0_share1_1 , x1x2x4_subscript0_share1_1 , x1x2x6_subscript0_share1_1 , x1x3x4_subscript0_share1_1 , x1x3x7_subscript0_share1_1 , x1x4x6_subscript0_share1_1 , x1x5x6_subscript0_share1_1 , x2x3x5_subscript0_share1_1 , x2x3x7_subscript0_share1_1 , x2x4x7_subscript0_share1_1 , x2x5x6_subscript0_share1_1 , x2x5x7_subscript0_share1_1 , x2x6x7_subscript0_share1_1 , x3x4x7_subscript0_share1_1 , x3x5x7_subscript0_share1_1 , x3x6x7_subscript0_share1_1 , x4x5x6_subscript0_share1_1 , x5x6x7_subscript0_share1_1 , x0x1x3_subscript0_share1_1 , x0x2x3_subscript0_share1_1 , x0x4x5_subscript0_share1_1 , x0x5x7_subscript0_share1_1 , x0x6x7_subscript0_share1_1 , x1x3x5_subscript0_share1_1 , x1x3x6_subscript0_share1_1 , x1x4x7_subscript0_share1_1 , x2x3x4_subscript0_share1_1 , x2x3x6_subscript0_share1_1 , x3x4x6_subscript0_share1_1 , x3x5x6_subscript0_share1_1 , x0x1x5_subscript0_share1_1 , x0x3x7_subscript0_share1_1 , x1x2x5_subscript0_share1_1 , x1x2x7_subscript0_share1_1 , x1x4x5_subscript0_share1_1 , x1x5x7_subscript0_share1_1 , x2x4x5_subscript0_share1_1 , x3x4x5_subscript0_share1_1 , x4x6x7_subscript0_share1_1 , x1x6x7_subscript0_share1_1 , x4x5x7_subscript0_share1_1 , x0x1x2_subscript0_share1_1 , x0x5x6_subscript0_share1_1 , x2x4x6_subscript0_share1_1 , x0x1x2x3_subscript0_share1_1 , x0x1x2x5_subscript0_share1_1 , x0x1x2x6_subscript0_share1_1 , x0x1x2x7_subscript0_share1_1 , x0x1x4x5_subscript0_share1_1 , x0x1x4x7_subscript0_share1_1 , x0x2x3x5_subscript0_share1_1 , x0x2x3x7_subscript0_share1_1 , x0x2x4x5_subscript0_share1_1 , x0x2x4x7_subscript0_share1_1 , x0x2x5x6_subscript0_share1_1 , x0x2x5x7_subscript0_share1_1 , x0x3x4x6_subscript0_share1_1 , x0x3x5x6_subscript0_share1_1 , x0x4x5x6_subscript0_share1_1 , x0x4x5x7_subscript0_share1_1 , x0x4x6x7_subscript0_share1_1 , x1x2x3x5_subscript0_share1_1 , x1x2x3x6_subscript0_share1_1 , x1x2x3x7_subscript0_share1_1 , x1x2x4x6_subscript0_share1_1 , x1x2x4x7_subscript0_share1_1 , x1x2x6x7_subscript0_share1_1 , x1x3x4x6_subscript0_share1_1 , x1x3x6x7_subscript0_share1_1 , x1x4x5x6_subscript0_share1_1 , x1x4x5x7_subscript0_share1_1 , x1x5x6x7_subscript0_share1_1 , x2x3x5x7_subscript0_share1_1 , x2x3x6x7_subscript0_share1_1 , x2x4x5x6_subscript0_share1_1 , x2x4x5x7_subscript0_share1_1 , x3x5x6x7_subscript0_share1_1 , x0x1x3x4_subscript0_share1_1 , x0x1x3x6_subscript0_share1_1 , x0x1x5x6_subscript0_share1_1 , x0x2x3x6_subscript0_share1_1 , x0x3x4x5_subscript0_share1_1 , x1x2x5x6_subscript0_share1_1 , x1x2x5x7_subscript0_share1_1 , x1x3x4x5_subscript0_share1_1 , x1x3x4x7_subscript0_share1_1 , x1x3x5x6_subscript0_share1_1 , x1x3x5x7_subscript0_share1_1 , x1x4x6x7_subscript0_share1_1 , x2x3x4x5_subscript0_share1_1 , x2x3x4x7_subscript0_share1_1 , x2x4x6x7_subscript0_share1_1 , x3x4x5x6_subscript0_share1_1 , x3x4x5x7_subscript0_share1_1 , x3x4x6x7_subscript0_share1_1 , x0x1x3x5_subscript0_share1_1 , x0x1x4x6_subscript0_share1_1 , x0x2x3x4_subscript0_share1_1 , x0x2x4x6_subscript0_share1_1 , x0x3x4x7_subscript0_share1_1 , x0x3x5x7_subscript0_share1_1 , x1x2x3x4_subscript0_share1_1 , x2x3x4x6_subscript0_share1_1 , x2x3x5x6_subscript0_share1_1 , x2x5x6x7_subscript0_share1_1 , x4x5x6x7_subscript0_share1_1 , x0x1x2x4_subscript0_share1_1 , x0x1x6x7_subscript0_share1_1 , x0x2x6x7_subscript0_share1_1 , x0x3x6x7_subscript0_share1_1 , x0x5x6x7_subscript0_share1_1 , x1x2x4x5_subscript0_share1_1 , x0x1x3x7_subscript0_share1_1 , x0x1x5x7_subscript0_share1_1 , x0x1x2x3x4_subscript0_share1_1 , x0x1x2x3x6_subscript0_share1_1 , x0x1x2x3x7_subscript0_share1_1 , x0x1x2x4x5_subscript0_share1_1 , x0x1x2x4x7_subscript0_share1_1 , x0x1x2x5x7_subscript0_share1_1 , x0x1x2x6x7_subscript0_share1_1 , x0x1x3x4x6_subscript0_share1_1 , x0x1x3x5x6_subscript0_share1_1 , x0x1x3x5x7_subscript0_share1_1 , x0x1x3x6x7_subscript0_share1_1 , x0x1x4x5x6_subscript0_share1_1 , x0x1x5x6x7_subscript0_share1_1 , x0x2x3x4x5_subscript0_share1_1 , x0x2x3x4x6_subscript0_share1_1 , x0x2x4x5x7_subscript0_share1_1 , x0x2x4x6x7_subscript0_share1_1 , x0x3x4x5x6_subscript0_share1_1 , x0x3x4x5x7_subscript0_share1_1 , x0x3x4x6x7_subscript0_share1_1 , x0x3x5x6x7_subscript0_share1_1 , x1x2x3x5x6_subscript0_share1_1 , x1x2x3x5x7_subscript0_share1_1 , x1x2x4x5x6_subscript0_share1_1 , x1x2x4x6x7_subscript0_share1_1 , x1x2x5x6x7_subscript0_share1_1 , x1x3x4x5x7_subscript0_share1_1 , x2x3x4x5x6_subscript0_share1_1 , x2x3x4x5x7_subscript0_share1_1 , x2x4x5x6x7_subscript0_share1_1 , x0x1x2x4x6_subscript0_share1_1 , x0x1x3x4x7_subscript0_share1_1 , x0x2x3x4x7_subscript0_share1_1 , x0x2x3x5x7_subscript0_share1_1 , x0x2x3x6x7_subscript0_share1_1 , x0x2x4x5x6_subscript0_share1_1 , x0x2x5x6x7_subscript0_share1_1 , x0x4x5x6x7_subscript0_share1_1 , x1x2x3x4x6_subscript0_share1_1 , x1x3x4x5x6_subscript0_share1_1 , x2x3x4x6x7_subscript0_share1_1 , x0x1x2x3x5_subscript0_share1_1 , x0x1x4x6x7_subscript0_share1_1 , x1x2x3x4x5_subscript0_share1_1 , x1x2x3x6x7_subscript0_share1_1 , x1x2x4x5x7_subscript0_share1_1 , x1x3x4x6x7_subscript0_share1_1 , x1x3x5x6x7_subscript0_share1_1 , x1x4x5x6x7_subscript0_share1_1 , x2x3x5x6x7_subscript0_share1_1 , x3x4x5x6x7_subscript0_share1_1 , x0x1x2x5x6_subscript0_share1_1 , x0x1x3x4x5_subscript0_share1_1 , x0x1x4x5x7_subscript0_share1_1 , x0x2x3x5x6_subscript0_share1_1 , x1x2x3x4x7_subscript0_share1_1 , x0x1x2x3x4x6_subscript0_share1_1 , x0x1x2x3x4x7_subscript0_share1_1 , x0x1x2x3x5x7_subscript0_share1_1 , x0x1x2x3x6x7_subscript0_share1_1 , x0x1x2x4x5x7_subscript0_share1_1 , x0x1x2x5x6x7_subscript0_share1_1 , x0x1x3x4x6x7_subscript0_share1_1 , x0x1x4x5x6x7_subscript0_share1_1 , x0x2x3x4x5x6_subscript0_share1_1 , x0x2x3x4x5x7_subscript0_share1_1 , x0x2x3x5x6x7_subscript0_share1_1 , x1x2x3x4x6x7_subscript0_share1_1 , x1x2x4x5x6x7_subscript0_share1_1 , x1x3x4x5x6x7_subscript0_share1_1 , x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x5x6_subscript0_share1_1 , x0x1x2x4x6x7_subscript0_share1_1 , x0x1x3x4x5x6_subscript0_share1_1 , x0x2x3x4x6x7_subscript0_share1_1 , x1x2x3x4x5x6_subscript0_share1_1 , x1x2x3x5x6x7_subscript0_share1_1 , x0x1x2x3x4x5_subscript0_share1_1 , x0x1x2x4x5x6_subscript0_share1_1 , x0x1x3x4x5x7_subscript0_share1_1 , x0x1x3x5x6x7_subscript0_share1_1 , x0x2x4x5x6x7_subscript0_share1_1 , x1x2x3x4x5x7_subscript0_share1_1 , x0x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x4x6x7_subscript0_share1_1 , x0x1x2x4x5x6x7_subscript0_share1_1 , x0x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x5x6x7_subscript0_share1_1 , x0x1x3x4x5x6x7_subscript0_share1_1 , x1x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x4x5x6_subscript0_share1_1 , x0x1x2x3x4x5x7_subscript0_share1_1 , x0_subscript0_share2_1 , x2_subscript0_share2_1 , x3_subscript0_share2_1 , x4_subscript0_share2_1 , x6_subscript0_share2_1 , x7_subscript0_share2_1 , x1_subscript0_share2_1 , x5_subscript0_share2_1 , x0x1_subscript0_share2_1 , x0x4_subscript0_share2_1 , x0x5_subscript0_share2_1 , x0x6_subscript0_share2_1 , x1x2_subscript0_share2_1 , x1x3_subscript0_share2_1 , x1x4_subscript0_share2_1 , x1x6_subscript0_share2_1 , x2x3_subscript0_share2_1 , x2x4_subscript0_share2_1 , x2x6_subscript0_share2_1 , x2x7_subscript0_share2_1 , x4x6_subscript0_share2_1 , x5x6_subscript0_share2_1 , x5x7_subscript0_share2_1 , x6x7_subscript0_share2_1 , x0x2_subscript0_share2_1 , x0x3_subscript0_share2_1 , x0x7_subscript0_share2_1 , x1x7_subscript0_share2_1 , x3x7_subscript0_share2_1 , x4x5_subscript0_share2_1 , x3x4_subscript0_share2_1 , x4x7_subscript0_share2_1 , x3x6_subscript0_share2_1 , x1x5_subscript0_share2_1 , x2x5_subscript0_share2_1 , x3x5_subscript0_share2_1 , x0x1x4_subscript0_share2_1 , x0x1x6_subscript0_share2_1 , x0x1x7_subscript0_share2_1 , x0x2x4_subscript0_share2_1 , x0x2x5_subscript0_share2_1 , x0x2x6_subscript0_share2_1 , x0x2x7_subscript0_share2_1 , x0x3x4_subscript0_share2_1 , x0x3x5_subscript0_share2_1 , x0x3x6_subscript0_share2_1 , x0x4x6_subscript0_share2_1 , x0x4x7_subscript0_share2_1 , x1x2x3_subscript0_share2_1 , x1x2x4_subscript0_share2_1 , x1x2x6_subscript0_share2_1 , x1x3x4_subscript0_share2_1 , x1x3x7_subscript0_share2_1 , x1x4x6_subscript0_share2_1 , x1x5x6_subscript0_share2_1 , x2x3x5_subscript0_share2_1 , x2x3x7_subscript0_share2_1 , x2x4x7_subscript0_share2_1 , x2x5x6_subscript0_share2_1 , x2x5x7_subscript0_share2_1 , x2x6x7_subscript0_share2_1 , x3x4x7_subscript0_share2_1 , x3x5x7_subscript0_share2_1 , x3x6x7_subscript0_share2_1 , x4x5x6_subscript0_share2_1 , x5x6x7_subscript0_share2_1 , x0x1x3_subscript0_share2_1 , x0x2x3_subscript0_share2_1 , x0x4x5_subscript0_share2_1 , x0x5x7_subscript0_share2_1 , x0x6x7_subscript0_share2_1 , x1x3x5_subscript0_share2_1 , x1x3x6_subscript0_share2_1 , x1x4x7_subscript0_share2_1 , x2x3x4_subscript0_share2_1 , x2x3x6_subscript0_share2_1 , x3x4x6_subscript0_share2_1 , x3x5x6_subscript0_share2_1 , x0x1x5_subscript0_share2_1 , x0x3x7_subscript0_share2_1 , x1x2x5_subscript0_share2_1 , x1x2x7_subscript0_share2_1 , x1x4x5_subscript0_share2_1 , x1x5x7_subscript0_share2_1 , x2x4x5_subscript0_share2_1 , x3x4x5_subscript0_share2_1 , x4x6x7_subscript0_share2_1 , x1x6x7_subscript0_share2_1 , x4x5x7_subscript0_share2_1 , x0x1x2_subscript0_share2_1 , x0x5x6_subscript0_share2_1 , x2x4x6_subscript0_share2_1 , x0x1x2x3_subscript0_share2_1 , x0x1x2x5_subscript0_share2_1 , x0x1x2x6_subscript0_share2_1 , x0x1x2x7_subscript0_share2_1 , x0x1x4x5_subscript0_share2_1 , x0x1x4x7_subscript0_share2_1 , x0x2x3x5_subscript0_share2_1 , x0x2x3x7_subscript0_share2_1 , x0x2x4x5_subscript0_share2_1 , x0x2x4x7_subscript0_share2_1 , x0x2x5x6_subscript0_share2_1 , x0x2x5x7_subscript0_share2_1 , x0x3x4x6_subscript0_share2_1 , x0x3x5x6_subscript0_share2_1 , x0x4x5x6_subscript0_share2_1 , x0x4x5x7_subscript0_share2_1 , x0x4x6x7_subscript0_share2_1 , x1x2x3x5_subscript0_share2_1 , x1x2x3x6_subscript0_share2_1 , x1x2x3x7_subscript0_share2_1 , x1x2x4x6_subscript0_share2_1 , x1x2x4x7_subscript0_share2_1 , x1x2x6x7_subscript0_share2_1 , x1x3x4x6_subscript0_share2_1 , x1x3x6x7_subscript0_share2_1 , x1x4x5x6_subscript0_share2_1 , x1x4x5x7_subscript0_share2_1 , x1x5x6x7_subscript0_share2_1 , x2x3x5x7_subscript0_share2_1 , x2x3x6x7_subscript0_share2_1 , x2x4x5x6_subscript0_share2_1 , x2x4x5x7_subscript0_share2_1 , x3x5x6x7_subscript0_share2_1 , x0x1x3x4_subscript0_share2_1 , x0x1x3x6_subscript0_share2_1 , x0x1x5x6_subscript0_share2_1 , x0x2x3x6_subscript0_share2_1 , x0x3x4x5_subscript0_share2_1 , x1x2x5x6_subscript0_share2_1 , x1x2x5x7_subscript0_share2_1 , x1x3x4x5_subscript0_share2_1 , x1x3x4x7_subscript0_share2_1 , x1x3x5x6_subscript0_share2_1 , x1x3x5x7_subscript0_share2_1 , x1x4x6x7_subscript0_share2_1 , x2x3x4x5_subscript0_share2_1 , x2x3x4x7_subscript0_share2_1 , x2x4x6x7_subscript0_share2_1 , x3x4x5x6_subscript0_share2_1 , x3x4x5x7_subscript0_share2_1 , x3x4x6x7_subscript0_share2_1 , x0x1x3x5_subscript0_share2_1 , x0x1x4x6_subscript0_share2_1 , x0x2x3x4_subscript0_share2_1 , x0x2x4x6_subscript0_share2_1 , x0x3x4x7_subscript0_share2_1 , x0x3x5x7_subscript0_share2_1 , x1x2x3x4_subscript0_share2_1 , x2x3x4x6_subscript0_share2_1 , x2x3x5x6_subscript0_share2_1 , x2x5x6x7_subscript0_share2_1 , x4x5x6x7_subscript0_share2_1 , x0x1x2x4_subscript0_share2_1 , x0x1x6x7_subscript0_share2_1 , x0x2x6x7_subscript0_share2_1 , x0x3x6x7_subscript0_share2_1 , x0x5x6x7_subscript0_share2_1 , x1x2x4x5_subscript0_share2_1 , x0x1x3x7_subscript0_share2_1 , x0x1x5x7_subscript0_share2_1 , x0x1x2x3x4_subscript0_share2_1 , x0x1x2x3x6_subscript0_share2_1 , x0x1x2x3x7_subscript0_share2_1 , x0x1x2x4x5_subscript0_share2_1 , x0x1x2x4x7_subscript0_share2_1 , x0x1x2x5x7_subscript0_share2_1 , x0x1x2x6x7_subscript0_share2_1 , x0x1x3x4x6_subscript0_share2_1 , x0x1x3x5x6_subscript0_share2_1 , x0x1x3x5x7_subscript0_share2_1 , x0x1x3x6x7_subscript0_share2_1 , x0x1x4x5x6_subscript0_share2_1 , x0x1x5x6x7_subscript0_share2_1 , x0x2x3x4x5_subscript0_share2_1 , x0x2x3x4x6_subscript0_share2_1 , x0x2x4x5x7_subscript0_share2_1 , x0x2x4x6x7_subscript0_share2_1 , x0x3x4x5x6_subscript0_share2_1 , x0x3x4x5x7_subscript0_share2_1 , x0x3x4x6x7_subscript0_share2_1 , x0x3x5x6x7_subscript0_share2_1 , x1x2x3x5x6_subscript0_share2_1 , x1x2x3x5x7_subscript0_share2_1 , x1x2x4x5x6_subscript0_share2_1 , x1x2x4x6x7_subscript0_share2_1 , x1x2x5x6x7_subscript0_share2_1 , x1x3x4x5x7_subscript0_share2_1 , x2x3x4x5x6_subscript0_share2_1 , x2x3x4x5x7_subscript0_share2_1 , x2x4x5x6x7_subscript0_share2_1 , x0x1x2x4x6_subscript0_share2_1 , x0x1x3x4x7_subscript0_share2_1 , x0x2x3x4x7_subscript0_share2_1 , x0x2x3x5x7_subscript0_share2_1 , x0x2x3x6x7_subscript0_share2_1 , x0x2x4x5x6_subscript0_share2_1 , x0x2x5x6x7_subscript0_share2_1 , x0x4x5x6x7_subscript0_share2_1 , x1x2x3x4x6_subscript0_share2_1 , x1x3x4x5x6_subscript0_share2_1 , x2x3x4x6x7_subscript0_share2_1 , x0x1x2x3x5_subscript0_share2_1 , x0x1x4x6x7_subscript0_share2_1 , x1x2x3x4x5_subscript0_share2_1 , x1x2x3x6x7_subscript0_share2_1 , x1x2x4x5x7_subscript0_share2_1 , x1x3x4x6x7_subscript0_share2_1 , x1x3x5x6x7_subscript0_share2_1 , x1x4x5x6x7_subscript0_share2_1 , x2x3x5x6x7_subscript0_share2_1 , x3x4x5x6x7_subscript0_share2_1 , x0x1x2x5x6_subscript0_share2_1 , x0x1x3x4x5_subscript0_share2_1 , x0x1x4x5x7_subscript0_share2_1 , x0x2x3x5x6_subscript0_share2_1 , x1x2x3x4x7_subscript0_share2_1 , x0x1x2x3x4x6_subscript0_share2_1 , x0x1x2x3x4x7_subscript0_share2_1 , x0x1x2x3x5x7_subscript0_share2_1 , x0x1x2x3x6x7_subscript0_share2_1 , x0x1x2x4x5x7_subscript0_share2_1 , x0x1x2x5x6x7_subscript0_share2_1 , x0x1x3x4x6x7_subscript0_share2_1 , x0x1x4x5x6x7_subscript0_share2_1 , x0x2x3x4x5x6_subscript0_share2_1 , x0x2x3x4x5x7_subscript0_share2_1 , x0x2x3x5x6x7_subscript0_share2_1 , x1x2x3x4x6x7_subscript0_share2_1 , x1x2x4x5x6x7_subscript0_share2_1 , x1x3x4x5x6x7_subscript0_share2_1 , x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x5x6_subscript0_share2_1 , x0x1x2x4x6x7_subscript0_share2_1 , x0x1x3x4x5x6_subscript0_share2_1 , x0x2x3x4x6x7_subscript0_share2_1 , x1x2x3x4x5x6_subscript0_share2_1 , x1x2x3x5x6x7_subscript0_share2_1 , x0x1x2x3x4x5_subscript0_share2_1 , x0x1x2x4x5x6_subscript0_share2_1 , x0x1x3x4x5x7_subscript0_share2_1 , x0x1x3x5x6x7_subscript0_share2_1 , x0x2x4x5x6x7_subscript0_share2_1 , x1x2x3x4x5x7_subscript0_share2_1 , x0x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x4x6x7_subscript0_share2_1 , x0x1x2x4x5x6x7_subscript0_share2_1 , x0x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x5x6x7_subscript0_share2_1 , x0x1x3x4x5x6x7_subscript0_share2_1 , x1x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x4x5x6_subscript0_share2_1 , x0x1x2x3x4x5x7_subscript0_share2_1 );
opt_AES_sbox_compute_subscript1 inst1( x0_subscript0_share1_reg , x2_subscript0_share1_reg , x3_subscript0_share1_reg , x4_subscript0_share1_reg , x6_subscript0_share1_reg , x7_subscript0_share1_reg , x1_subscript0_share1_reg , x5_subscript0_share1_reg , x0x1_subscript0_share1_reg , x0x4_subscript0_share1_reg , x0x5_subscript0_share1_reg , x0x6_subscript0_share1_reg , x1x2_subscript0_share1_reg , x1x3_subscript0_share1_reg , x1x4_subscript0_share1_reg , x1x6_subscript0_share1_reg , x2x3_subscript0_share1_reg , x2x4_subscript0_share1_reg , x2x6_subscript0_share1_reg , x2x7_subscript0_share1_reg , x4x6_subscript0_share1_reg , x5x6_subscript0_share1_reg , x5x7_subscript0_share1_reg , x6x7_subscript0_share1_reg , x0x2_subscript0_share1_reg , x0x3_subscript0_share1_reg , x0x7_subscript0_share1_reg , x1x7_subscript0_share1_reg , x3x7_subscript0_share1_reg , x4x5_subscript0_share1_reg , x3x4_subscript0_share1_reg , x4x7_subscript0_share1_reg , x3x6_subscript0_share1_reg , x1x5_subscript0_share1_reg , x2x5_subscript0_share1_reg , x3x5_subscript0_share1_reg , x0x1x4_subscript0_share1_reg , x0x1x6_subscript0_share1_reg , x0x1x7_subscript0_share1_reg , x0x2x4_subscript0_share1_reg , x0x2x5_subscript0_share1_reg , x0x2x6_subscript0_share1_reg , x0x2x7_subscript0_share1_reg , x0x3x4_subscript0_share1_reg , x0x3x5_subscript0_share1_reg , x0x3x6_subscript0_share1_reg , x0x4x6_subscript0_share1_reg , x0x4x7_subscript0_share1_reg , x1x2x3_subscript0_share1_reg , x1x2x4_subscript0_share1_reg , x1x2x6_subscript0_share1_reg , x1x3x4_subscript0_share1_reg , x1x3x7_subscript0_share1_reg , x1x4x6_subscript0_share1_reg , x1x5x6_subscript0_share1_reg , x2x3x5_subscript0_share1_reg , x2x3x7_subscript0_share1_reg , x2x4x7_subscript0_share1_reg , x2x5x6_subscript0_share1_reg , x2x5x7_subscript0_share1_reg , x2x6x7_subscript0_share1_reg , x3x4x7_subscript0_share1_reg , x3x5x7_subscript0_share1_reg , x3x6x7_subscript0_share1_reg , x4x5x6_subscript0_share1_reg , x5x6x7_subscript0_share1_reg , x0x1x3_subscript0_share1_reg , x0x2x3_subscript0_share1_reg , x0x4x5_subscript0_share1_reg , x0x5x7_subscript0_share1_reg , x0x6x7_subscript0_share1_reg , x1x3x5_subscript0_share1_reg , x1x3x6_subscript0_share1_reg , x1x4x7_subscript0_share1_reg , x2x3x4_subscript0_share1_reg , x2x3x6_subscript0_share1_reg , x3x4x6_subscript0_share1_reg , x3x5x6_subscript0_share1_reg , x0x1x5_subscript0_share1_reg , x0x3x7_subscript0_share1_reg , x1x2x5_subscript0_share1_reg , x1x2x7_subscript0_share1_reg , x1x4x5_subscript0_share1_reg , x1x5x7_subscript0_share1_reg , x2x4x5_subscript0_share1_reg , x3x4x5_subscript0_share1_reg , x4x6x7_subscript0_share1_reg , x1x6x7_subscript0_share1_reg , x4x5x7_subscript0_share1_reg , x0x1x2_subscript0_share1_reg , x0x5x6_subscript0_share1_reg , x2x4x6_subscript0_share1_reg , x0x1x2x3_subscript0_share1_reg , x0x1x2x5_subscript0_share1_reg , x0x1x2x6_subscript0_share1_reg , x0x1x2x7_subscript0_share1_reg , x0x1x4x5_subscript0_share1_reg , x0x1x4x7_subscript0_share1_reg , x0x2x3x5_subscript0_share1_reg , x0x2x3x7_subscript0_share1_reg , x0x2x4x5_subscript0_share1_reg , x0x2x4x7_subscript0_share1_reg , x0x2x5x6_subscript0_share1_reg , x0x2x5x7_subscript0_share1_reg , x0x3x4x6_subscript0_share1_reg , x0x3x5x6_subscript0_share1_reg , x0x4x5x6_subscript0_share1_reg , x0x4x5x7_subscript0_share1_reg , x0x4x6x7_subscript0_share1_reg , x1x2x3x5_subscript0_share1_reg , x1x2x3x6_subscript0_share1_reg , x1x2x3x7_subscript0_share1_reg , x1x2x4x6_subscript0_share1_reg , x1x2x4x7_subscript0_share1_reg , x1x2x6x7_subscript0_share1_reg , x1x3x4x6_subscript0_share1_reg , x1x3x6x7_subscript0_share1_reg , x1x4x5x6_subscript0_share1_reg , x1x4x5x7_subscript0_share1_reg , x1x5x6x7_subscript0_share1_reg , x2x3x5x7_subscript0_share1_reg , x2x3x6x7_subscript0_share1_reg , x2x4x5x6_subscript0_share1_reg , x2x4x5x7_subscript0_share1_reg , x3x5x6x7_subscript0_share1_reg , x0x1x3x4_subscript0_share1_reg , x0x1x3x6_subscript0_share1_reg , x0x1x5x6_subscript0_share1_reg , x0x2x3x6_subscript0_share1_reg , x0x3x4x5_subscript0_share1_reg , x1x2x5x6_subscript0_share1_reg , x1x2x5x7_subscript0_share1_reg , x1x3x4x5_subscript0_share1_reg , x1x3x4x7_subscript0_share1_reg , x1x3x5x6_subscript0_share1_reg , x1x3x5x7_subscript0_share1_reg , x1x4x6x7_subscript0_share1_reg , x2x3x4x5_subscript0_share1_reg , x2x3x4x7_subscript0_share1_reg , x2x4x6x7_subscript0_share1_reg , x3x4x5x6_subscript0_share1_reg , x3x4x5x7_subscript0_share1_reg , x3x4x6x7_subscript0_share1_reg , x0x1x3x5_subscript0_share1_reg , x0x1x4x6_subscript0_share1_reg , x0x2x3x4_subscript0_share1_reg , x0x2x4x6_subscript0_share1_reg , x0x3x4x7_subscript0_share1_reg , x0x3x5x7_subscript0_share1_reg , x1x2x3x4_subscript0_share1_reg , x2x3x4x6_subscript0_share1_reg , x2x3x5x6_subscript0_share1_reg , x2x5x6x7_subscript0_share1_reg , x4x5x6x7_subscript0_share1_reg , x0x1x2x4_subscript0_share1_reg , x0x1x6x7_subscript0_share1_reg , x0x2x6x7_subscript0_share1_reg , x0x3x6x7_subscript0_share1_reg , x0x5x6x7_subscript0_share1_reg , x1x2x4x5_subscript0_share1_reg , x0x1x3x7_subscript0_share1_reg , x0x1x5x7_subscript0_share1_reg , x0x1x2x3x4_subscript0_share1_reg , x0x1x2x3x6_subscript0_share1_reg , x0x1x2x3x7_subscript0_share1_reg , x0x1x2x4x5_subscript0_share1_reg , x0x1x2x4x7_subscript0_share1_reg , x0x1x2x5x7_subscript0_share1_reg , x0x1x2x6x7_subscript0_share1_reg , x0x1x3x4x6_subscript0_share1_reg , x0x1x3x5x6_subscript0_share1_reg , x0x1x3x5x7_subscript0_share1_reg , x0x1x3x6x7_subscript0_share1_reg , x0x1x4x5x6_subscript0_share1_reg , x0x1x5x6x7_subscript0_share1_reg , x0x2x3x4x5_subscript0_share1_reg , x0x2x3x4x6_subscript0_share1_reg , x0x2x4x5x7_subscript0_share1_reg , x0x2x4x6x7_subscript0_share1_reg , x0x3x4x5x6_subscript0_share1_reg , x0x3x4x5x7_subscript0_share1_reg , x0x3x4x6x7_subscript0_share1_reg , x0x3x5x6x7_subscript0_share1_reg , x1x2x3x5x6_subscript0_share1_reg , x1x2x3x5x7_subscript0_share1_reg , x1x2x4x5x6_subscript0_share1_reg , x1x2x4x6x7_subscript0_share1_reg , x1x2x5x6x7_subscript0_share1_reg , x1x3x4x5x7_subscript0_share1_reg , x2x3x4x5x6_subscript0_share1_reg , x2x3x4x5x7_subscript0_share1_reg , x2x4x5x6x7_subscript0_share1_reg , x0x1x2x4x6_subscript0_share1_reg , x0x1x3x4x7_subscript0_share1_reg , x0x2x3x4x7_subscript0_share1_reg , x0x2x3x5x7_subscript0_share1_reg , x0x2x3x6x7_subscript0_share1_reg , x0x2x4x5x6_subscript0_share1_reg , x0x2x5x6x7_subscript0_share1_reg , x0x4x5x6x7_subscript0_share1_reg , x1x2x3x4x6_subscript0_share1_reg , x1x3x4x5x6_subscript0_share1_reg , x2x3x4x6x7_subscript0_share1_reg , x0x1x2x3x5_subscript0_share1_reg , x0x1x4x6x7_subscript0_share1_reg , x1x2x3x4x5_subscript0_share1_reg , x1x2x3x6x7_subscript0_share1_reg , x1x2x4x5x7_subscript0_share1_reg , x1x3x4x6x7_subscript0_share1_reg , x1x3x5x6x7_subscript0_share1_reg , x1x4x5x6x7_subscript0_share1_reg , x2x3x5x6x7_subscript0_share1_reg , x3x4x5x6x7_subscript0_share1_reg , x0x1x2x5x6_subscript0_share1_reg , x0x1x3x4x5_subscript0_share1_reg , x0x1x4x5x7_subscript0_share1_reg , x0x2x3x5x6_subscript0_share1_reg , x1x2x3x4x7_subscript0_share1_reg , x0x1x2x3x4x6_subscript0_share1_reg , x0x1x2x3x4x7_subscript0_share1_reg , x0x1x2x3x5x7_subscript0_share1_reg , x0x1x2x3x6x7_subscript0_share1_reg , x0x1x2x4x5x7_subscript0_share1_reg , x0x1x2x5x6x7_subscript0_share1_reg , x0x1x3x4x6x7_subscript0_share1_reg , x0x1x4x5x6x7_subscript0_share1_reg , x0x2x3x4x5x6_subscript0_share1_reg , x0x2x3x4x5x7_subscript0_share1_reg , x0x2x3x5x6x7_subscript0_share1_reg , x1x2x3x4x6x7_subscript0_share1_reg , x1x2x4x5x6x7_subscript0_share1_reg , x1x3x4x5x6x7_subscript0_share1_reg , x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x5x6_subscript0_share1_reg , x0x1x2x4x6x7_subscript0_share1_reg , x0x1x3x4x5x6_subscript0_share1_reg , x0x2x3x4x6x7_subscript0_share1_reg , x1x2x3x4x5x6_subscript0_share1_reg , x1x2x3x5x6x7_subscript0_share1_reg , x0x1x2x3x4x5_subscript0_share1_reg , x0x1x2x4x5x6_subscript0_share1_reg , x0x1x3x4x5x7_subscript0_share1_reg , x0x1x3x5x6x7_subscript0_share1_reg , x0x2x4x5x6x7_subscript0_share1_reg , x1x2x3x4x5x7_subscript0_share1_reg , x0x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x4x6x7_subscript0_share1_reg , x0x1x2x4x5x6x7_subscript0_share1_reg , x0x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x5x6x7_subscript0_share1_reg , x0x1x3x4x5x6x7_subscript0_share1_reg , x1x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x4x5x6_subscript0_share1_reg , x0x1x2x3x4x5x7_subscript0_share1_reg , x0_subscript0_share2_reg , x2_subscript0_share2_reg , x3_subscript0_share2_reg , x4_subscript0_share2_reg , x6_subscript0_share2_reg , x7_subscript0_share2_reg , x1_subscript0_share2_reg , x5_subscript0_share2_reg , x0x1_subscript0_share2_reg , x0x4_subscript0_share2_reg , x0x5_subscript0_share2_reg , x0x6_subscript0_share2_reg , x1x2_subscript0_share2_reg , x1x3_subscript0_share2_reg , x1x4_subscript0_share2_reg , x1x6_subscript0_share2_reg , x2x3_subscript0_share2_reg , x2x4_subscript0_share2_reg , x2x6_subscript0_share2_reg , x2x7_subscript0_share2_reg , x4x6_subscript0_share2_reg , x5x6_subscript0_share2_reg , x5x7_subscript0_share2_reg , x6x7_subscript0_share2_reg , x0x2_subscript0_share2_reg , x0x3_subscript0_share2_reg , x0x7_subscript0_share2_reg , x1x7_subscript0_share2_reg , x3x7_subscript0_share2_reg , x4x5_subscript0_share2_reg , x3x4_subscript0_share2_reg , x4x7_subscript0_share2_reg , x3x6_subscript0_share2_reg , x1x5_subscript0_share2_reg , x2x5_subscript0_share2_reg , x3x5_subscript0_share2_reg , x0x1x4_subscript0_share2_reg , x0x1x6_subscript0_share2_reg , x0x1x7_subscript0_share2_reg , x0x2x4_subscript0_share2_reg , x0x2x5_subscript0_share2_reg , x0x2x6_subscript0_share2_reg , x0x2x7_subscript0_share2_reg , x0x3x4_subscript0_share2_reg , x0x3x5_subscript0_share2_reg , x0x3x6_subscript0_share2_reg , x0x4x6_subscript0_share2_reg , x0x4x7_subscript0_share2_reg , x1x2x3_subscript0_share2_reg , x1x2x4_subscript0_share2_reg , x1x2x6_subscript0_share2_reg , x1x3x4_subscript0_share2_reg , x1x3x7_subscript0_share2_reg , x1x4x6_subscript0_share2_reg , x1x5x6_subscript0_share2_reg , x2x3x5_subscript0_share2_reg , x2x3x7_subscript0_share2_reg , x2x4x7_subscript0_share2_reg , x2x5x6_subscript0_share2_reg , x2x5x7_subscript0_share2_reg , x2x6x7_subscript0_share2_reg , x3x4x7_subscript0_share2_reg , x3x5x7_subscript0_share2_reg , x3x6x7_subscript0_share2_reg , x4x5x6_subscript0_share2_reg , x5x6x7_subscript0_share2_reg , x0x1x3_subscript0_share2_reg , x0x2x3_subscript0_share2_reg , x0x4x5_subscript0_share2_reg , x0x5x7_subscript0_share2_reg , x0x6x7_subscript0_share2_reg , x1x3x5_subscript0_share2_reg , x1x3x6_subscript0_share2_reg , x1x4x7_subscript0_share2_reg , x2x3x4_subscript0_share2_reg , x2x3x6_subscript0_share2_reg , x3x4x6_subscript0_share2_reg , x3x5x6_subscript0_share2_reg , x0x1x5_subscript0_share2_reg , x0x3x7_subscript0_share2_reg , x1x2x5_subscript0_share2_reg , x1x2x7_subscript0_share2_reg , x1x4x5_subscript0_share2_reg , x1x5x7_subscript0_share2_reg , x2x4x5_subscript0_share2_reg , x3x4x5_subscript0_share2_reg , x4x6x7_subscript0_share2_reg , x1x6x7_subscript0_share2_reg , x4x5x7_subscript0_share2_reg , x0x1x2_subscript0_share2_reg , x0x5x6_subscript0_share2_reg , x2x4x6_subscript0_share2_reg , x0x1x2x3_subscript0_share2_reg , x0x1x2x5_subscript0_share2_reg , x0x1x2x6_subscript0_share2_reg , x0x1x2x7_subscript0_share2_reg , x0x1x4x5_subscript0_share2_reg , x0x1x4x7_subscript0_share2_reg , x0x2x3x5_subscript0_share2_reg , x0x2x3x7_subscript0_share2_reg , x0x2x4x5_subscript0_share2_reg , x0x2x4x7_subscript0_share2_reg , x0x2x5x6_subscript0_share2_reg , x0x2x5x7_subscript0_share2_reg , x0x3x4x6_subscript0_share2_reg , x0x3x5x6_subscript0_share2_reg , x0x4x5x6_subscript0_share2_reg , x0x4x5x7_subscript0_share2_reg , x0x4x6x7_subscript0_share2_reg , x1x2x3x5_subscript0_share2_reg , x1x2x3x6_subscript0_share2_reg , x1x2x3x7_subscript0_share2_reg , x1x2x4x6_subscript0_share2_reg , x1x2x4x7_subscript0_share2_reg , x1x2x6x7_subscript0_share2_reg , x1x3x4x6_subscript0_share2_reg , x1x3x6x7_subscript0_share2_reg , x1x4x5x6_subscript0_share2_reg , x1x4x5x7_subscript0_share2_reg , x1x5x6x7_subscript0_share2_reg , x2x3x5x7_subscript0_share2_reg , x2x3x6x7_subscript0_share2_reg , x2x4x5x6_subscript0_share2_reg , x2x4x5x7_subscript0_share2_reg , x3x5x6x7_subscript0_share2_reg , x0x1x3x4_subscript0_share2_reg , x0x1x3x6_subscript0_share2_reg , x0x1x5x6_subscript0_share2_reg , x0x2x3x6_subscript0_share2_reg , x0x3x4x5_subscript0_share2_reg , x1x2x5x6_subscript0_share2_reg , x1x2x5x7_subscript0_share2_reg , x1x3x4x5_subscript0_share2_reg , x1x3x4x7_subscript0_share2_reg , x1x3x5x6_subscript0_share2_reg , x1x3x5x7_subscript0_share2_reg , x1x4x6x7_subscript0_share2_reg , x2x3x4x5_subscript0_share2_reg , x2x3x4x7_subscript0_share2_reg , x2x4x6x7_subscript0_share2_reg , x3x4x5x6_subscript0_share2_reg , x3x4x5x7_subscript0_share2_reg , x3x4x6x7_subscript0_share2_reg , x0x1x3x5_subscript0_share2_reg , x0x1x4x6_subscript0_share2_reg , x0x2x3x4_subscript0_share2_reg , x0x2x4x6_subscript0_share2_reg , x0x3x4x7_subscript0_share2_reg , x0x3x5x7_subscript0_share2_reg , x1x2x3x4_subscript0_share2_reg , x2x3x4x6_subscript0_share2_reg , x2x3x5x6_subscript0_share2_reg , x2x5x6x7_subscript0_share2_reg , x4x5x6x7_subscript0_share2_reg , x0x1x2x4_subscript0_share2_reg , x0x1x6x7_subscript0_share2_reg , x0x2x6x7_subscript0_share2_reg , x0x3x6x7_subscript0_share2_reg , x0x5x6x7_subscript0_share2_reg , x1x2x4x5_subscript0_share2_reg , x0x1x3x7_subscript0_share2_reg , x0x1x5x7_subscript0_share2_reg , x0x1x2x3x4_subscript0_share2_reg , x0x1x2x3x6_subscript0_share2_reg , x0x1x2x3x7_subscript0_share2_reg , x0x1x2x4x5_subscript0_share2_reg , x0x1x2x4x7_subscript0_share2_reg , x0x1x2x5x7_subscript0_share2_reg , x0x1x2x6x7_subscript0_share2_reg , x0x1x3x4x6_subscript0_share2_reg , x0x1x3x5x6_subscript0_share2_reg , x0x1x3x5x7_subscript0_share2_reg , x0x1x3x6x7_subscript0_share2_reg , x0x1x4x5x6_subscript0_share2_reg , x0x1x5x6x7_subscript0_share2_reg , x0x2x3x4x5_subscript0_share2_reg , x0x2x3x4x6_subscript0_share2_reg , x0x2x4x5x7_subscript0_share2_reg , x0x2x4x6x7_subscript0_share2_reg , x0x3x4x5x6_subscript0_share2_reg , x0x3x4x5x7_subscript0_share2_reg , x0x3x4x6x7_subscript0_share2_reg , x0x3x5x6x7_subscript0_share2_reg , x1x2x3x5x6_subscript0_share2_reg , x1x2x3x5x7_subscript0_share2_reg , x1x2x4x5x6_subscript0_share2_reg , x1x2x4x6x7_subscript0_share2_reg , x1x2x5x6x7_subscript0_share2_reg , x1x3x4x5x7_subscript0_share2_reg , x2x3x4x5x6_subscript0_share2_reg , x2x3x4x5x7_subscript0_share2_reg , x2x4x5x6x7_subscript0_share2_reg , x0x1x2x4x6_subscript0_share2_reg , x0x1x3x4x7_subscript0_share2_reg , x0x2x3x4x7_subscript0_share2_reg , x0x2x3x5x7_subscript0_share2_reg , x0x2x3x6x7_subscript0_share2_reg , x0x2x4x5x6_subscript0_share2_reg , x0x2x5x6x7_subscript0_share2_reg , x0x4x5x6x7_subscript0_share2_reg , x1x2x3x4x6_subscript0_share2_reg , x1x3x4x5x6_subscript0_share2_reg , x2x3x4x6x7_subscript0_share2_reg , x0x1x2x3x5_subscript0_share2_reg , x0x1x4x6x7_subscript0_share2_reg , x1x2x3x4x5_subscript0_share2_reg , x1x2x3x6x7_subscript0_share2_reg , x1x2x4x5x7_subscript0_share2_reg , x1x3x4x6x7_subscript0_share2_reg , x1x3x5x6x7_subscript0_share2_reg , x1x4x5x6x7_subscript0_share2_reg , x2x3x5x6x7_subscript0_share2_reg , x3x4x5x6x7_subscript0_share2_reg , x0x1x2x5x6_subscript0_share2_reg , x0x1x3x4x5_subscript0_share2_reg , x0x1x4x5x7_subscript0_share2_reg , x0x2x3x5x6_subscript0_share2_reg , x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x4x6_subscript0_share2_reg , x0x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x5x7_subscript0_share2_reg , x0x1x2x3x6x7_subscript0_share2_reg , x0x1x2x4x5x7_subscript0_share2_reg , x0x1x2x5x6x7_subscript0_share2_reg , x0x1x3x4x6x7_subscript0_share2_reg , x0x1x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6_subscript0_share2_reg , x0x2x3x4x5x7_subscript0_share2_reg , x0x2x3x5x6x7_subscript0_share2_reg , x1x2x3x4x6x7_subscript0_share2_reg , x1x2x4x5x6x7_subscript0_share2_reg , x1x3x4x5x6x7_subscript0_share2_reg , x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6_subscript0_share2_reg , x0x1x2x4x6x7_subscript0_share2_reg , x0x1x3x4x5x6_subscript0_share2_reg , x0x2x3x4x6x7_subscript0_share2_reg , x1x2x3x4x5x6_subscript0_share2_reg , x1x2x3x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5_subscript0_share2_reg , x0x1x2x4x5x6_subscript0_share2_reg , x0x1x3x4x5x7_subscript0_share2_reg , x0x1x3x5x6x7_subscript0_share2_reg , x0x2x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x7_subscript0_share2_reg , x0x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x6x7_subscript0_share2_reg , x0x1x2x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6x7_subscript0_share2_reg , x0x1x3x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5x6_subscript0_share2_reg , x0x1x2x3x4x5x7_subscript0_share2_reg ,x0_share2_reg , x1_share2_reg , x2_share2_reg , x3_share2_reg , x4_share2_reg , x5_share2_reg , x6_share2_reg , x7_share2_reg ,    sbox_out1_share1, sbox_out2_share1, sbox_out3_share1, sbox_out4_share1, sbox_out5_share1, sbox_out6_share1, sbox_out7_share1, sbox_out8_share1 ,     sbox_out1_share2, sbox_out2_share2, sbox_out3_share2, sbox_out4_share2, sbox_out5_share2, sbox_out6_share2, sbox_out7_share2, sbox_out8_share2  );


always@(posedge clk) begin
                
        x0_share2_reg <= sbox_input_share2[0] ^ rand_composable_bit[0] ;
        x1_share2_reg <= sbox_input_share2[1] ^ rand_composable_bit[1] ;
        x2_share2_reg <= sbox_input_share2[2] ^ rand_composable_bit[2] ;
        x3_share2_reg <= sbox_input_share2[3] ^ rand_composable_bit[3] ;
        x4_share2_reg <= sbox_input_share2[4] ^ rand_composable_bit[4] ;
        x5_share2_reg <= sbox_input_share2[5] ^ rand_composable_bit[5] ;
        x6_share2_reg <= sbox_input_share2[6] ^ rand_composable_bit[6] ;
        x7_share2_reg <= sbox_input_share2[7] ^ rand_composable_bit[7] ;

        x0_subscript0_share1_reg <= x0_subscript0_share1_1 ; 
        x0_subscript0_share2_reg <= x0_subscript0_share2_1 ; 
        x2_subscript0_share1_reg <= x2_subscript0_share1_1 ; 
        x2_subscript0_share2_reg <= x2_subscript0_share2_1 ; 
        x3_subscript0_share1_reg <= x3_subscript0_share1_1 ; 
        x3_subscript0_share2_reg <= x3_subscript0_share2_1 ; 
        x4_subscript0_share1_reg <= x4_subscript0_share1_1 ; 
        x4_subscript0_share2_reg <= x4_subscript0_share2_1 ; 
        x6_subscript0_share1_reg <= x6_subscript0_share1_1 ; 
        x6_subscript0_share2_reg <= x6_subscript0_share2_1 ; 
        x7_subscript0_share1_reg <= x7_subscript0_share1_1 ; 
        x7_subscript0_share2_reg <= x7_subscript0_share2_1 ; 
        x1_subscript0_share1_reg <= x1_subscript0_share1_1 ; 
        x1_subscript0_share2_reg <= x1_subscript0_share2_1 ; 
        x5_subscript0_share1_reg <= x5_subscript0_share1_1 ; 
        x5_subscript0_share2_reg <= x5_subscript0_share2_1 ; 
        x0x1_subscript0_share1_reg <= x0x1_subscript0_share1_1 ; 
        x0x1_subscript0_share2_reg <= x0x1_subscript0_share2_1 ; 
        x0x4_subscript0_share1_reg <= x0x4_subscript0_share1_1 ; 
        x0x4_subscript0_share2_reg <= x0x4_subscript0_share2_1 ; 
        x0x5_subscript0_share1_reg <= x0x5_subscript0_share1_1 ; 
        x0x5_subscript0_share2_reg <= x0x5_subscript0_share2_1 ; 
        x0x6_subscript0_share1_reg <= x0x6_subscript0_share1_1 ; 
        x0x6_subscript0_share2_reg <= x0x6_subscript0_share2_1 ; 
        x1x2_subscript0_share1_reg <= x1x2_subscript0_share1_1 ; 
        x1x2_subscript0_share2_reg <= x1x2_subscript0_share2_1 ; 
        x1x3_subscript0_share1_reg <= x1x3_subscript0_share1_1 ; 
        x1x3_subscript0_share2_reg <= x1x3_subscript0_share2_1 ; 
        x1x4_subscript0_share1_reg <= x1x4_subscript0_share1_1 ; 
        x1x4_subscript0_share2_reg <= x1x4_subscript0_share2_1 ; 
        x1x6_subscript0_share1_reg <= x1x6_subscript0_share1_1 ; 
        x1x6_subscript0_share2_reg <= x1x6_subscript0_share2_1 ; 
        x2x3_subscript0_share1_reg <= x2x3_subscript0_share1_1 ; 
        x2x3_subscript0_share2_reg <= x2x3_subscript0_share2_1 ; 
        x2x4_subscript0_share1_reg <= x2x4_subscript0_share1_1 ; 
        x2x4_subscript0_share2_reg <= x2x4_subscript0_share2_1 ; 
        x2x6_subscript0_share1_reg <= x2x6_subscript0_share1_1 ; 
        x2x6_subscript0_share2_reg <= x2x6_subscript0_share2_1 ; 
        x2x7_subscript0_share1_reg <= x2x7_subscript0_share1_1 ; 
        x2x7_subscript0_share2_reg <= x2x7_subscript0_share2_1 ; 
        x4x6_subscript0_share1_reg <= x4x6_subscript0_share1_1 ; 
        x4x6_subscript0_share2_reg <= x4x6_subscript0_share2_1 ; 
        x5x6_subscript0_share1_reg <= x5x6_subscript0_share1_1 ; 
        x5x6_subscript0_share2_reg <= x5x6_subscript0_share2_1 ; 
        x5x7_subscript0_share1_reg <= x5x7_subscript0_share1_1 ; 
        x5x7_subscript0_share2_reg <= x5x7_subscript0_share2_1 ; 
        x6x7_subscript0_share1_reg <= x6x7_subscript0_share1_1 ; 
        x6x7_subscript0_share2_reg <= x6x7_subscript0_share2_1 ; 
        x0x2_subscript0_share1_reg <= x0x2_subscript0_share1_1 ; 
        x0x2_subscript0_share2_reg <= x0x2_subscript0_share2_1 ; 
        x0x3_subscript0_share1_reg <= x0x3_subscript0_share1_1 ; 
        x0x3_subscript0_share2_reg <= x0x3_subscript0_share2_1 ; 
        x0x7_subscript0_share1_reg <= x0x7_subscript0_share1_1 ; 
        x0x7_subscript0_share2_reg <= x0x7_subscript0_share2_1 ; 
        x1x7_subscript0_share1_reg <= x1x7_subscript0_share1_1 ; 
        x1x7_subscript0_share2_reg <= x1x7_subscript0_share2_1 ; 
        x3x7_subscript0_share1_reg <= x3x7_subscript0_share1_1 ; 
        x3x7_subscript0_share2_reg <= x3x7_subscript0_share2_1 ; 
        x4x5_subscript0_share1_reg <= x4x5_subscript0_share1_1 ; 
        x4x5_subscript0_share2_reg <= x4x5_subscript0_share2_1 ; 
        x3x4_subscript0_share1_reg <= x3x4_subscript0_share1_1 ; 
        x3x4_subscript0_share2_reg <= x3x4_subscript0_share2_1 ; 
        x4x7_subscript0_share1_reg <= x4x7_subscript0_share1_1 ; 
        x4x7_subscript0_share2_reg <= x4x7_subscript0_share2_1 ; 
        x3x6_subscript0_share1_reg <= x3x6_subscript0_share1_1 ; 
        x3x6_subscript0_share2_reg <= x3x6_subscript0_share2_1 ; 
        x1x5_subscript0_share1_reg <= x1x5_subscript0_share1_1 ; 
        x1x5_subscript0_share2_reg <= x1x5_subscript0_share2_1 ; 
        x2x5_subscript0_share1_reg <= x2x5_subscript0_share1_1 ; 
        x2x5_subscript0_share2_reg <= x2x5_subscript0_share2_1 ; 
        x3x5_subscript0_share1_reg <= x3x5_subscript0_share1_1 ; 
        x3x5_subscript0_share2_reg <= x3x5_subscript0_share2_1 ; 
        x0x1x4_subscript0_share1_reg <= x0x1x4_subscript0_share1_1 ; 
        x0x1x4_subscript0_share2_reg <= x0x1x4_subscript0_share2_1 ; 
        x0x1x6_subscript0_share1_reg <= x0x1x6_subscript0_share1_1 ; 
        x0x1x6_subscript0_share2_reg <= x0x1x6_subscript0_share2_1 ; 
        x0x1x7_subscript0_share1_reg <= x0x1x7_subscript0_share1_1 ; 
        x0x1x7_subscript0_share2_reg <= x0x1x7_subscript0_share2_1 ; 
        x0x2x4_subscript0_share1_reg <= x0x2x4_subscript0_share1_1 ; 
        x0x2x4_subscript0_share2_reg <= x0x2x4_subscript0_share2_1 ; 
        x0x2x5_subscript0_share1_reg <= x0x2x5_subscript0_share1_1 ; 
        x0x2x5_subscript0_share2_reg <= x0x2x5_subscript0_share2_1 ; 
        x0x2x6_subscript0_share1_reg <= x0x2x6_subscript0_share1_1 ; 
        x0x2x6_subscript0_share2_reg <= x0x2x6_subscript0_share2_1 ; 
        x0x2x7_subscript0_share1_reg <= x0x2x7_subscript0_share1_1 ; 
        x0x2x7_subscript0_share2_reg <= x0x2x7_subscript0_share2_1 ; 
        x0x3x4_subscript0_share1_reg <= x0x3x4_subscript0_share1_1 ; 
        x0x3x4_subscript0_share2_reg <= x0x3x4_subscript0_share2_1 ; 
        x0x3x5_subscript0_share1_reg <= x0x3x5_subscript0_share1_1 ; 
        x0x3x5_subscript0_share2_reg <= x0x3x5_subscript0_share2_1 ; 
        x0x3x6_subscript0_share1_reg <= x0x3x6_subscript0_share1_1 ; 
        x0x3x6_subscript0_share2_reg <= x0x3x6_subscript0_share2_1 ; 
        x0x4x6_subscript0_share1_reg <= x0x4x6_subscript0_share1_1 ; 
        x0x4x6_subscript0_share2_reg <= x0x4x6_subscript0_share2_1 ; 
        x0x4x7_subscript0_share1_reg <= x0x4x7_subscript0_share1_1 ; 
        x0x4x7_subscript0_share2_reg <= x0x4x7_subscript0_share2_1 ; 
        x1x2x3_subscript0_share1_reg <= x1x2x3_subscript0_share1_1 ; 
        x1x2x3_subscript0_share2_reg <= x1x2x3_subscript0_share2_1 ; 
        x1x2x4_subscript0_share1_reg <= x1x2x4_subscript0_share1_1 ; 
        x1x2x4_subscript0_share2_reg <= x1x2x4_subscript0_share2_1 ; 
        x1x2x6_subscript0_share1_reg <= x1x2x6_subscript0_share1_1 ; 
        x1x2x6_subscript0_share2_reg <= x1x2x6_subscript0_share2_1 ; 
        x1x3x4_subscript0_share1_reg <= x1x3x4_subscript0_share1_1 ; 
        x1x3x4_subscript0_share2_reg <= x1x3x4_subscript0_share2_1 ; 
        x1x3x7_subscript0_share1_reg <= x1x3x7_subscript0_share1_1 ; 
        x1x3x7_subscript0_share2_reg <= x1x3x7_subscript0_share2_1 ; 
        x1x4x6_subscript0_share1_reg <= x1x4x6_subscript0_share1_1 ; 
        x1x4x6_subscript0_share2_reg <= x1x4x6_subscript0_share2_1 ; 
        x1x5x6_subscript0_share1_reg <= x1x5x6_subscript0_share1_1 ; 
        x1x5x6_subscript0_share2_reg <= x1x5x6_subscript0_share2_1 ; 
        x2x3x5_subscript0_share1_reg <= x2x3x5_subscript0_share1_1 ; 
        x2x3x5_subscript0_share2_reg <= x2x3x5_subscript0_share2_1 ; 
        x2x3x7_subscript0_share1_reg <= x2x3x7_subscript0_share1_1 ; 
        x2x3x7_subscript0_share2_reg <= x2x3x7_subscript0_share2_1 ; 
        x2x4x7_subscript0_share1_reg <= x2x4x7_subscript0_share1_1 ; 
        x2x4x7_subscript0_share2_reg <= x2x4x7_subscript0_share2_1 ; 
        x2x5x6_subscript0_share1_reg <= x2x5x6_subscript0_share1_1 ; 
        x2x5x6_subscript0_share2_reg <= x2x5x6_subscript0_share2_1 ; 
        x2x5x7_subscript0_share1_reg <= x2x5x7_subscript0_share1_1 ; 
        x2x5x7_subscript0_share2_reg <= x2x5x7_subscript0_share2_1 ; 
        x2x6x7_subscript0_share1_reg <= x2x6x7_subscript0_share1_1 ; 
        x2x6x7_subscript0_share2_reg <= x2x6x7_subscript0_share2_1 ; 
        x3x4x7_subscript0_share1_reg <= x3x4x7_subscript0_share1_1 ; 
        x3x4x7_subscript0_share2_reg <= x3x4x7_subscript0_share2_1 ; 
        x3x5x7_subscript0_share1_reg <= x3x5x7_subscript0_share1_1 ; 
        x3x5x7_subscript0_share2_reg <= x3x5x7_subscript0_share2_1 ; 
        x3x6x7_subscript0_share1_reg <= x3x6x7_subscript0_share1_1 ; 
        x3x6x7_subscript0_share2_reg <= x3x6x7_subscript0_share2_1 ; 
        x4x5x6_subscript0_share1_reg <= x4x5x6_subscript0_share1_1 ; 
        x4x5x6_subscript0_share2_reg <= x4x5x6_subscript0_share2_1 ; 
        x5x6x7_subscript0_share1_reg <= x5x6x7_subscript0_share1_1 ; 
        x5x6x7_subscript0_share2_reg <= x5x6x7_subscript0_share2_1 ; 
        x0x1x3_subscript0_share1_reg <= x0x1x3_subscript0_share1_1 ; 
        x0x1x3_subscript0_share2_reg <= x0x1x3_subscript0_share2_1 ; 
        x0x2x3_subscript0_share1_reg <= x0x2x3_subscript0_share1_1 ; 
        x0x2x3_subscript0_share2_reg <= x0x2x3_subscript0_share2_1 ; 
        x0x4x5_subscript0_share1_reg <= x0x4x5_subscript0_share1_1 ; 
        x0x4x5_subscript0_share2_reg <= x0x4x5_subscript0_share2_1 ; 
        x0x5x7_subscript0_share1_reg <= x0x5x7_subscript0_share1_1 ; 
        x0x5x7_subscript0_share2_reg <= x0x5x7_subscript0_share2_1 ; 
        x0x6x7_subscript0_share1_reg <= x0x6x7_subscript0_share1_1 ; 
        x0x6x7_subscript0_share2_reg <= x0x6x7_subscript0_share2_1 ; 
        x1x3x5_subscript0_share1_reg <= x1x3x5_subscript0_share1_1 ; 
        x1x3x5_subscript0_share2_reg <= x1x3x5_subscript0_share2_1 ; 
        x1x3x6_subscript0_share1_reg <= x1x3x6_subscript0_share1_1 ; 
        x1x3x6_subscript0_share2_reg <= x1x3x6_subscript0_share2_1 ; 
        x1x4x7_subscript0_share1_reg <= x1x4x7_subscript0_share1_1 ; 
        x1x4x7_subscript0_share2_reg <= x1x4x7_subscript0_share2_1 ; 
        x2x3x4_subscript0_share1_reg <= x2x3x4_subscript0_share1_1 ; 
        x2x3x4_subscript0_share2_reg <= x2x3x4_subscript0_share2_1 ; 
        x2x3x6_subscript0_share1_reg <= x2x3x6_subscript0_share1_1 ; 
        x2x3x6_subscript0_share2_reg <= x2x3x6_subscript0_share2_1 ; 
        x3x4x6_subscript0_share1_reg <= x3x4x6_subscript0_share1_1 ; 
        x3x4x6_subscript0_share2_reg <= x3x4x6_subscript0_share2_1 ; 
        x3x5x6_subscript0_share1_reg <= x3x5x6_subscript0_share1_1 ; 
        x3x5x6_subscript0_share2_reg <= x3x5x6_subscript0_share2_1 ; 
        x0x1x5_subscript0_share1_reg <= x0x1x5_subscript0_share1_1 ; 
        x0x1x5_subscript0_share2_reg <= x0x1x5_subscript0_share2_1 ; 
        x0x3x7_subscript0_share1_reg <= x0x3x7_subscript0_share1_1 ; 
        x0x3x7_subscript0_share2_reg <= x0x3x7_subscript0_share2_1 ; 
        x1x2x5_subscript0_share1_reg <= x1x2x5_subscript0_share1_1 ; 
        x1x2x5_subscript0_share2_reg <= x1x2x5_subscript0_share2_1 ; 
        x1x2x7_subscript0_share1_reg <= x1x2x7_subscript0_share1_1 ; 
        x1x2x7_subscript0_share2_reg <= x1x2x7_subscript0_share2_1 ; 
        x1x4x5_subscript0_share1_reg <= x1x4x5_subscript0_share1_1 ; 
        x1x4x5_subscript0_share2_reg <= x1x4x5_subscript0_share2_1 ; 
        x1x5x7_subscript0_share1_reg <= x1x5x7_subscript0_share1_1 ; 
        x1x5x7_subscript0_share2_reg <= x1x5x7_subscript0_share2_1 ; 
        x2x4x5_subscript0_share1_reg <= x2x4x5_subscript0_share1_1 ; 
        x2x4x5_subscript0_share2_reg <= x2x4x5_subscript0_share2_1 ; 
        x3x4x5_subscript0_share1_reg <= x3x4x5_subscript0_share1_1 ; 
        x3x4x5_subscript0_share2_reg <= x3x4x5_subscript0_share2_1 ; 
        x4x6x7_subscript0_share1_reg <= x4x6x7_subscript0_share1_1 ; 
        x4x6x7_subscript0_share2_reg <= x4x6x7_subscript0_share2_1 ; 
        x1x6x7_subscript0_share1_reg <= x1x6x7_subscript0_share1_1 ; 
        x1x6x7_subscript0_share2_reg <= x1x6x7_subscript0_share2_1 ; 
        x4x5x7_subscript0_share1_reg <= x4x5x7_subscript0_share1_1 ; 
        x4x5x7_subscript0_share2_reg <= x4x5x7_subscript0_share2_1 ; 
        x0x1x2_subscript0_share1_reg <= x0x1x2_subscript0_share1_1 ; 
        x0x1x2_subscript0_share2_reg <= x0x1x2_subscript0_share2_1 ; 
        x0x5x6_subscript0_share1_reg <= x0x5x6_subscript0_share1_1 ; 
        x0x5x6_subscript0_share2_reg <= x0x5x6_subscript0_share2_1 ; 
        x2x4x6_subscript0_share1_reg <= x2x4x6_subscript0_share1_1 ; 
        x2x4x6_subscript0_share2_reg <= x2x4x6_subscript0_share2_1 ; 
        x0x1x2x3_subscript0_share1_reg <= x0x1x2x3_subscript0_share1_1 ; 
        x0x1x2x3_subscript0_share2_reg <= x0x1x2x3_subscript0_share2_1 ; 
        x0x1x2x5_subscript0_share1_reg <= x0x1x2x5_subscript0_share1_1 ; 
        x0x1x2x5_subscript0_share2_reg <= x0x1x2x5_subscript0_share2_1 ; 
        x0x1x2x6_subscript0_share1_reg <= x0x1x2x6_subscript0_share1_1 ; 
        x0x1x2x6_subscript0_share2_reg <= x0x1x2x6_subscript0_share2_1 ; 
        x0x1x2x7_subscript0_share1_reg <= x0x1x2x7_subscript0_share1_1 ; 
        x0x1x2x7_subscript0_share2_reg <= x0x1x2x7_subscript0_share2_1 ; 
        x0x1x4x5_subscript0_share1_reg <= x0x1x4x5_subscript0_share1_1 ; 
        x0x1x4x5_subscript0_share2_reg <= x0x1x4x5_subscript0_share2_1 ; 
        x0x1x4x7_subscript0_share1_reg <= x0x1x4x7_subscript0_share1_1 ; 
        x0x1x4x7_subscript0_share2_reg <= x0x1x4x7_subscript0_share2_1 ; 
        x0x2x3x5_subscript0_share1_reg <= x0x2x3x5_subscript0_share1_1 ; 
        x0x2x3x5_subscript0_share2_reg <= x0x2x3x5_subscript0_share2_1 ; 
        x0x2x3x7_subscript0_share1_reg <= x0x2x3x7_subscript0_share1_1 ; 
        x0x2x3x7_subscript0_share2_reg <= x0x2x3x7_subscript0_share2_1 ; 
        x0x2x4x5_subscript0_share1_reg <= x0x2x4x5_subscript0_share1_1 ; 
        x0x2x4x5_subscript0_share2_reg <= x0x2x4x5_subscript0_share2_1 ; 
        x0x2x4x7_subscript0_share1_reg <= x0x2x4x7_subscript0_share1_1 ; 
        x0x2x4x7_subscript0_share2_reg <= x0x2x4x7_subscript0_share2_1 ; 
        x0x2x5x6_subscript0_share1_reg <= x0x2x5x6_subscript0_share1_1 ; 
        x0x2x5x6_subscript0_share2_reg <= x0x2x5x6_subscript0_share2_1 ; 
        x0x2x5x7_subscript0_share1_reg <= x0x2x5x7_subscript0_share1_1 ; 
        x0x2x5x7_subscript0_share2_reg <= x0x2x5x7_subscript0_share2_1 ; 
        x0x3x4x6_subscript0_share1_reg <= x0x3x4x6_subscript0_share1_1 ; 
        x0x3x4x6_subscript0_share2_reg <= x0x3x4x6_subscript0_share2_1 ; 
        x0x3x5x6_subscript0_share1_reg <= x0x3x5x6_subscript0_share1_1 ; 
        x0x3x5x6_subscript0_share2_reg <= x0x3x5x6_subscript0_share2_1 ; 
        x0x4x5x6_subscript0_share1_reg <= x0x4x5x6_subscript0_share1_1 ; 
        x0x4x5x6_subscript0_share2_reg <= x0x4x5x6_subscript0_share2_1 ; 
        x0x4x5x7_subscript0_share1_reg <= x0x4x5x7_subscript0_share1_1 ; 
        x0x4x5x7_subscript0_share2_reg <= x0x4x5x7_subscript0_share2_1 ; 
        x0x4x6x7_subscript0_share1_reg <= x0x4x6x7_subscript0_share1_1 ; 
        x0x4x6x7_subscript0_share2_reg <= x0x4x6x7_subscript0_share2_1 ; 
        x1x2x3x5_subscript0_share1_reg <= x1x2x3x5_subscript0_share1_1 ; 
        x1x2x3x5_subscript0_share2_reg <= x1x2x3x5_subscript0_share2_1 ; 
        x1x2x3x6_subscript0_share1_reg <= x1x2x3x6_subscript0_share1_1 ; 
        x1x2x3x6_subscript0_share2_reg <= x1x2x3x6_subscript0_share2_1 ; 
        x1x2x3x7_subscript0_share1_reg <= x1x2x3x7_subscript0_share1_1 ; 
        x1x2x3x7_subscript0_share2_reg <= x1x2x3x7_subscript0_share2_1 ; 
        x1x2x4x6_subscript0_share1_reg <= x1x2x4x6_subscript0_share1_1 ; 
        x1x2x4x6_subscript0_share2_reg <= x1x2x4x6_subscript0_share2_1 ; 
        x1x2x4x7_subscript0_share1_reg <= x1x2x4x7_subscript0_share1_1 ; 
        x1x2x4x7_subscript0_share2_reg <= x1x2x4x7_subscript0_share2_1 ; 
        x1x2x6x7_subscript0_share1_reg <= x1x2x6x7_subscript0_share1_1 ; 
        x1x2x6x7_subscript0_share2_reg <= x1x2x6x7_subscript0_share2_1 ; 
        x1x3x4x6_subscript0_share1_reg <= x1x3x4x6_subscript0_share1_1 ; 
        x1x3x4x6_subscript0_share2_reg <= x1x3x4x6_subscript0_share2_1 ; 
        x1x3x6x7_subscript0_share1_reg <= x1x3x6x7_subscript0_share1_1 ; 
        x1x3x6x7_subscript0_share2_reg <= x1x3x6x7_subscript0_share2_1 ; 
        x1x4x5x6_subscript0_share1_reg <= x1x4x5x6_subscript0_share1_1 ; 
        x1x4x5x6_subscript0_share2_reg <= x1x4x5x6_subscript0_share2_1 ; 
        x1x4x5x7_subscript0_share1_reg <= x1x4x5x7_subscript0_share1_1 ; 
        x1x4x5x7_subscript0_share2_reg <= x1x4x5x7_subscript0_share2_1 ; 
        x1x5x6x7_subscript0_share1_reg <= x1x5x6x7_subscript0_share1_1 ; 
        x1x5x6x7_subscript0_share2_reg <= x1x5x6x7_subscript0_share2_1 ; 
        x2x3x5x7_subscript0_share1_reg <= x2x3x5x7_subscript0_share1_1 ; 
        x2x3x5x7_subscript0_share2_reg <= x2x3x5x7_subscript0_share2_1 ; 
        x2x3x6x7_subscript0_share1_reg <= x2x3x6x7_subscript0_share1_1 ; 
        x2x3x6x7_subscript0_share2_reg <= x2x3x6x7_subscript0_share2_1 ; 
        x2x4x5x6_subscript0_share1_reg <= x2x4x5x6_subscript0_share1_1 ; 
        x2x4x5x6_subscript0_share2_reg <= x2x4x5x6_subscript0_share2_1 ; 
        x2x4x5x7_subscript0_share1_reg <= x2x4x5x7_subscript0_share1_1 ; 
        x2x4x5x7_subscript0_share2_reg <= x2x4x5x7_subscript0_share2_1 ; 
        x3x5x6x7_subscript0_share1_reg <= x3x5x6x7_subscript0_share1_1 ; 
        x3x5x6x7_subscript0_share2_reg <= x3x5x6x7_subscript0_share2_1 ; 
        x0x1x3x4_subscript0_share1_reg <= x0x1x3x4_subscript0_share1_1 ; 
        x0x1x3x4_subscript0_share2_reg <= x0x1x3x4_subscript0_share2_1 ; 
        x0x1x3x6_subscript0_share1_reg <= x0x1x3x6_subscript0_share1_1 ; 
        x0x1x3x6_subscript0_share2_reg <= x0x1x3x6_subscript0_share2_1 ; 
        x0x1x5x6_subscript0_share1_reg <= x0x1x5x6_subscript0_share1_1 ; 
        x0x1x5x6_subscript0_share2_reg <= x0x1x5x6_subscript0_share2_1 ; 
        x0x2x3x6_subscript0_share1_reg <= x0x2x3x6_subscript0_share1_1 ; 
        x0x2x3x6_subscript0_share2_reg <= x0x2x3x6_subscript0_share2_1 ; 
        x0x3x4x5_subscript0_share1_reg <= x0x3x4x5_subscript0_share1_1 ; 
        x0x3x4x5_subscript0_share2_reg <= x0x3x4x5_subscript0_share2_1 ; 
        x1x2x5x6_subscript0_share1_reg <= x1x2x5x6_subscript0_share1_1 ; 
        x1x2x5x6_subscript0_share2_reg <= x1x2x5x6_subscript0_share2_1 ; 
        x1x2x5x7_subscript0_share1_reg <= x1x2x5x7_subscript0_share1_1 ; 
        x1x2x5x7_subscript0_share2_reg <= x1x2x5x7_subscript0_share2_1 ; 
        x1x3x4x5_subscript0_share1_reg <= x1x3x4x5_subscript0_share1_1 ; 
        x1x3x4x5_subscript0_share2_reg <= x1x3x4x5_subscript0_share2_1 ; 
        x1x3x4x7_subscript0_share1_reg <= x1x3x4x7_subscript0_share1_1 ; 
        x1x3x4x7_subscript0_share2_reg <= x1x3x4x7_subscript0_share2_1 ; 
        x1x3x5x6_subscript0_share1_reg <= x1x3x5x6_subscript0_share1_1 ; 
        x1x3x5x6_subscript0_share2_reg <= x1x3x5x6_subscript0_share2_1 ; 
        x1x3x5x7_subscript0_share1_reg <= x1x3x5x7_subscript0_share1_1 ; 
        x1x3x5x7_subscript0_share2_reg <= x1x3x5x7_subscript0_share2_1 ; 
        x1x4x6x7_subscript0_share1_reg <= x1x4x6x7_subscript0_share1_1 ; 
        x1x4x6x7_subscript0_share2_reg <= x1x4x6x7_subscript0_share2_1 ; 
        x2x3x4x5_subscript0_share1_reg <= x2x3x4x5_subscript0_share1_1 ; 
        x2x3x4x5_subscript0_share2_reg <= x2x3x4x5_subscript0_share2_1 ; 
        x2x3x4x7_subscript0_share1_reg <= x2x3x4x7_subscript0_share1_1 ; 
        x2x3x4x7_subscript0_share2_reg <= x2x3x4x7_subscript0_share2_1 ; 
        x2x4x6x7_subscript0_share1_reg <= x2x4x6x7_subscript0_share1_1 ; 
        x2x4x6x7_subscript0_share2_reg <= x2x4x6x7_subscript0_share2_1 ; 
        x3x4x5x6_subscript0_share1_reg <= x3x4x5x6_subscript0_share1_1 ; 
        x3x4x5x6_subscript0_share2_reg <= x3x4x5x6_subscript0_share2_1 ; 
        x3x4x5x7_subscript0_share1_reg <= x3x4x5x7_subscript0_share1_1 ; 
        x3x4x5x7_subscript0_share2_reg <= x3x4x5x7_subscript0_share2_1 ; 
        x3x4x6x7_subscript0_share1_reg <= x3x4x6x7_subscript0_share1_1 ; 
        x3x4x6x7_subscript0_share2_reg <= x3x4x6x7_subscript0_share2_1 ; 
        x0x1x3x5_subscript0_share1_reg <= x0x1x3x5_subscript0_share1_1 ; 
        x0x1x3x5_subscript0_share2_reg <= x0x1x3x5_subscript0_share2_1 ; 
        x0x1x4x6_subscript0_share1_reg <= x0x1x4x6_subscript0_share1_1 ; 
        x0x1x4x6_subscript0_share2_reg <= x0x1x4x6_subscript0_share2_1 ; 
        x0x2x3x4_subscript0_share1_reg <= x0x2x3x4_subscript0_share1_1 ; 
        x0x2x3x4_subscript0_share2_reg <= x0x2x3x4_subscript0_share2_1 ; 
        x0x2x4x6_subscript0_share1_reg <= x0x2x4x6_subscript0_share1_1 ; 
        x0x2x4x6_subscript0_share2_reg <= x0x2x4x6_subscript0_share2_1 ; 
        x0x3x4x7_subscript0_share1_reg <= x0x3x4x7_subscript0_share1_1 ; 
        x0x3x4x7_subscript0_share2_reg <= x0x3x4x7_subscript0_share2_1 ; 
        x0x3x5x7_subscript0_share1_reg <= x0x3x5x7_subscript0_share1_1 ; 
        x0x3x5x7_subscript0_share2_reg <= x0x3x5x7_subscript0_share2_1 ; 
        x1x2x3x4_subscript0_share1_reg <= x1x2x3x4_subscript0_share1_1 ; 
        x1x2x3x4_subscript0_share2_reg <= x1x2x3x4_subscript0_share2_1 ; 
        x2x3x4x6_subscript0_share1_reg <= x2x3x4x6_subscript0_share1_1 ; 
        x2x3x4x6_subscript0_share2_reg <= x2x3x4x6_subscript0_share2_1 ; 
        x2x3x5x6_subscript0_share1_reg <= x2x3x5x6_subscript0_share1_1 ; 
        x2x3x5x6_subscript0_share2_reg <= x2x3x5x6_subscript0_share2_1 ; 
        x2x5x6x7_subscript0_share1_reg <= x2x5x6x7_subscript0_share1_1 ; 
        x2x5x6x7_subscript0_share2_reg <= x2x5x6x7_subscript0_share2_1 ; 
        x4x5x6x7_subscript0_share1_reg <= x4x5x6x7_subscript0_share1_1 ; 
        x4x5x6x7_subscript0_share2_reg <= x4x5x6x7_subscript0_share2_1 ; 
        x0x1x2x4_subscript0_share1_reg <= x0x1x2x4_subscript0_share1_1 ; 
        x0x1x2x4_subscript0_share2_reg <= x0x1x2x4_subscript0_share2_1 ; 
        x0x1x6x7_subscript0_share1_reg <= x0x1x6x7_subscript0_share1_1 ; 
        x0x1x6x7_subscript0_share2_reg <= x0x1x6x7_subscript0_share2_1 ; 
        x0x2x6x7_subscript0_share1_reg <= x0x2x6x7_subscript0_share1_1 ; 
        x0x2x6x7_subscript0_share2_reg <= x0x2x6x7_subscript0_share2_1 ; 
        x0x3x6x7_subscript0_share1_reg <= x0x3x6x7_subscript0_share1_1 ; 
        x0x3x6x7_subscript0_share2_reg <= x0x3x6x7_subscript0_share2_1 ; 
        x0x5x6x7_subscript0_share1_reg <= x0x5x6x7_subscript0_share1_1 ; 
        x0x5x6x7_subscript0_share2_reg <= x0x5x6x7_subscript0_share2_1 ; 
        x1x2x4x5_subscript0_share1_reg <= x1x2x4x5_subscript0_share1_1 ; 
        x1x2x4x5_subscript0_share2_reg <= x1x2x4x5_subscript0_share2_1 ; 
        x0x1x3x7_subscript0_share1_reg <= x0x1x3x7_subscript0_share1_1 ; 
        x0x1x3x7_subscript0_share2_reg <= x0x1x3x7_subscript0_share2_1 ; 
        x0x1x5x7_subscript0_share1_reg <= x0x1x5x7_subscript0_share1_1 ; 
        x0x1x5x7_subscript0_share2_reg <= x0x1x5x7_subscript0_share2_1 ; 
        x0x1x2x3x4_subscript0_share1_reg <= x0x1x2x3x4_subscript0_share1_1 ; 
        x0x1x2x3x4_subscript0_share2_reg <= x0x1x2x3x4_subscript0_share2_1 ; 
        x0x1x2x3x6_subscript0_share1_reg <= x0x1x2x3x6_subscript0_share1_1 ; 
        x0x1x2x3x6_subscript0_share2_reg <= x0x1x2x3x6_subscript0_share2_1 ; 
        x0x1x2x3x7_subscript0_share1_reg <= x0x1x2x3x7_subscript0_share1_1 ; 
        x0x1x2x3x7_subscript0_share2_reg <= x0x1x2x3x7_subscript0_share2_1 ; 
        x0x1x2x4x5_subscript0_share1_reg <= x0x1x2x4x5_subscript0_share1_1 ; 
        x0x1x2x4x5_subscript0_share2_reg <= x0x1x2x4x5_subscript0_share2_1 ; 
        x0x1x2x4x7_subscript0_share1_reg <= x0x1x2x4x7_subscript0_share1_1 ; 
        x0x1x2x4x7_subscript0_share2_reg <= x0x1x2x4x7_subscript0_share2_1 ; 
        x0x1x2x5x7_subscript0_share1_reg <= x0x1x2x5x7_subscript0_share1_1 ; 
        x0x1x2x5x7_subscript0_share2_reg <= x0x1x2x5x7_subscript0_share2_1 ; 
        x0x1x2x6x7_subscript0_share1_reg <= x0x1x2x6x7_subscript0_share1_1 ; 
        x0x1x2x6x7_subscript0_share2_reg <= x0x1x2x6x7_subscript0_share2_1 ; 
        x0x1x3x4x6_subscript0_share1_reg <= x0x1x3x4x6_subscript0_share1_1 ; 
        x0x1x3x4x6_subscript0_share2_reg <= x0x1x3x4x6_subscript0_share2_1 ; 
        x0x1x3x5x6_subscript0_share1_reg <= x0x1x3x5x6_subscript0_share1_1 ; 
        x0x1x3x5x6_subscript0_share2_reg <= x0x1x3x5x6_subscript0_share2_1 ; 
        x0x1x3x5x7_subscript0_share1_reg <= x0x1x3x5x7_subscript0_share1_1 ; 
        x0x1x3x5x7_subscript0_share2_reg <= x0x1x3x5x7_subscript0_share2_1 ; 
        x0x1x3x6x7_subscript0_share1_reg <= x0x1x3x6x7_subscript0_share1_1 ; 
        x0x1x3x6x7_subscript0_share2_reg <= x0x1x3x6x7_subscript0_share2_1 ; 
        x0x1x4x5x6_subscript0_share1_reg <= x0x1x4x5x6_subscript0_share1_1 ; 
        x0x1x4x5x6_subscript0_share2_reg <= x0x1x4x5x6_subscript0_share2_1 ; 
        x0x1x5x6x7_subscript0_share1_reg <= x0x1x5x6x7_subscript0_share1_1 ; 
        x0x1x5x6x7_subscript0_share2_reg <= x0x1x5x6x7_subscript0_share2_1 ; 
        x0x2x3x4x5_subscript0_share1_reg <= x0x2x3x4x5_subscript0_share1_1 ; 
        x0x2x3x4x5_subscript0_share2_reg <= x0x2x3x4x5_subscript0_share2_1 ; 
        x0x2x3x4x6_subscript0_share1_reg <= x0x2x3x4x6_subscript0_share1_1 ; 
        x0x2x3x4x6_subscript0_share2_reg <= x0x2x3x4x6_subscript0_share2_1 ; 
        x0x2x4x5x7_subscript0_share1_reg <= x0x2x4x5x7_subscript0_share1_1 ; 
        x0x2x4x5x7_subscript0_share2_reg <= x0x2x4x5x7_subscript0_share2_1 ; 
        x0x2x4x6x7_subscript0_share1_reg <= x0x2x4x6x7_subscript0_share1_1 ; 
        x0x2x4x6x7_subscript0_share2_reg <= x0x2x4x6x7_subscript0_share2_1 ; 
        x0x3x4x5x6_subscript0_share1_reg <= x0x3x4x5x6_subscript0_share1_1 ; 
        x0x3x4x5x6_subscript0_share2_reg <= x0x3x4x5x6_subscript0_share2_1 ; 
        x0x3x4x5x7_subscript0_share1_reg <= x0x3x4x5x7_subscript0_share1_1 ; 
        x0x3x4x5x7_subscript0_share2_reg <= x0x3x4x5x7_subscript0_share2_1 ; 
        x0x3x4x6x7_subscript0_share1_reg <= x0x3x4x6x7_subscript0_share1_1 ; 
        x0x3x4x6x7_subscript0_share2_reg <= x0x3x4x6x7_subscript0_share2_1 ; 
        x0x3x5x6x7_subscript0_share1_reg <= x0x3x5x6x7_subscript0_share1_1 ; 
        x0x3x5x6x7_subscript0_share2_reg <= x0x3x5x6x7_subscript0_share2_1 ; 
        x1x2x3x5x6_subscript0_share1_reg <= x1x2x3x5x6_subscript0_share1_1 ; 
        x1x2x3x5x6_subscript0_share2_reg <= x1x2x3x5x6_subscript0_share2_1 ; 
        x1x2x3x5x7_subscript0_share1_reg <= x1x2x3x5x7_subscript0_share1_1 ; 
        x1x2x3x5x7_subscript0_share2_reg <= x1x2x3x5x7_subscript0_share2_1 ; 
        x1x2x4x5x6_subscript0_share1_reg <= x1x2x4x5x6_subscript0_share1_1 ; 
        x1x2x4x5x6_subscript0_share2_reg <= x1x2x4x5x6_subscript0_share2_1 ; 
        x1x2x4x6x7_subscript0_share1_reg <= x1x2x4x6x7_subscript0_share1_1 ; 
        x1x2x4x6x7_subscript0_share2_reg <= x1x2x4x6x7_subscript0_share2_1 ; 
        x1x2x5x6x7_subscript0_share1_reg <= x1x2x5x6x7_subscript0_share1_1 ; 
        x1x2x5x6x7_subscript0_share2_reg <= x1x2x5x6x7_subscript0_share2_1 ; 
        x1x3x4x5x7_subscript0_share1_reg <= x1x3x4x5x7_subscript0_share1_1 ; 
        x1x3x4x5x7_subscript0_share2_reg <= x1x3x4x5x7_subscript0_share2_1 ; 
        x2x3x4x5x6_subscript0_share1_reg <= x2x3x4x5x6_subscript0_share1_1 ; 
        x2x3x4x5x6_subscript0_share2_reg <= x2x3x4x5x6_subscript0_share2_1 ; 
        x2x3x4x5x7_subscript0_share1_reg <= x2x3x4x5x7_subscript0_share1_1 ; 
        x2x3x4x5x7_subscript0_share2_reg <= x2x3x4x5x7_subscript0_share2_1 ; 
        x2x4x5x6x7_subscript0_share1_reg <= x2x4x5x6x7_subscript0_share1_1 ; 
        x2x4x5x6x7_subscript0_share2_reg <= x2x4x5x6x7_subscript0_share2_1 ; 
        x0x1x2x4x6_subscript0_share1_reg <= x0x1x2x4x6_subscript0_share1_1 ; 
        x0x1x2x4x6_subscript0_share2_reg <= x0x1x2x4x6_subscript0_share2_1 ; 
        x0x1x3x4x7_subscript0_share1_reg <= x0x1x3x4x7_subscript0_share1_1 ; 
        x0x1x3x4x7_subscript0_share2_reg <= x0x1x3x4x7_subscript0_share2_1 ; 
        x0x2x3x4x7_subscript0_share1_reg <= x0x2x3x4x7_subscript0_share1_1 ; 
        x0x2x3x4x7_subscript0_share2_reg <= x0x2x3x4x7_subscript0_share2_1 ; 
        x0x2x3x5x7_subscript0_share1_reg <= x0x2x3x5x7_subscript0_share1_1 ; 
        x0x2x3x5x7_subscript0_share2_reg <= x0x2x3x5x7_subscript0_share2_1 ; 
        x0x2x3x6x7_subscript0_share1_reg <= x0x2x3x6x7_subscript0_share1_1 ; 
        x0x2x3x6x7_subscript0_share2_reg <= x0x2x3x6x7_subscript0_share2_1 ; 
        x0x2x4x5x6_subscript0_share1_reg <= x0x2x4x5x6_subscript0_share1_1 ; 
        x0x2x4x5x6_subscript0_share2_reg <= x0x2x4x5x6_subscript0_share2_1 ; 
        x0x2x5x6x7_subscript0_share1_reg <= x0x2x5x6x7_subscript0_share1_1 ; 
        x0x2x5x6x7_subscript0_share2_reg <= x0x2x5x6x7_subscript0_share2_1 ; 
        x0x4x5x6x7_subscript0_share1_reg <= x0x4x5x6x7_subscript0_share1_1 ; 
        x0x4x5x6x7_subscript0_share2_reg <= x0x4x5x6x7_subscript0_share2_1 ; 
        x1x2x3x4x6_subscript0_share1_reg <= x1x2x3x4x6_subscript0_share1_1 ; 
        x1x2x3x4x6_subscript0_share2_reg <= x1x2x3x4x6_subscript0_share2_1 ; 
        x1x3x4x5x6_subscript0_share1_reg <= x1x3x4x5x6_subscript0_share1_1 ; 
        x1x3x4x5x6_subscript0_share2_reg <= x1x3x4x5x6_subscript0_share2_1 ; 
        x2x3x4x6x7_subscript0_share1_reg <= x2x3x4x6x7_subscript0_share1_1 ; 
        x2x3x4x6x7_subscript0_share2_reg <= x2x3x4x6x7_subscript0_share2_1 ; 
        x0x1x2x3x5_subscript0_share1_reg <= x0x1x2x3x5_subscript0_share1_1 ; 
        x0x1x2x3x5_subscript0_share2_reg <= x0x1x2x3x5_subscript0_share2_1 ; 
        x0x1x4x6x7_subscript0_share1_reg <= x0x1x4x6x7_subscript0_share1_1 ; 
        x0x1x4x6x7_subscript0_share2_reg <= x0x1x4x6x7_subscript0_share2_1 ; 
        x1x2x3x4x5_subscript0_share1_reg <= x1x2x3x4x5_subscript0_share1_1 ; 
        x1x2x3x4x5_subscript0_share2_reg <= x1x2x3x4x5_subscript0_share2_1 ; 
        x1x2x3x6x7_subscript0_share1_reg <= x1x2x3x6x7_subscript0_share1_1 ; 
        x1x2x3x6x7_subscript0_share2_reg <= x1x2x3x6x7_subscript0_share2_1 ; 
        x1x2x4x5x7_subscript0_share1_reg <= x1x2x4x5x7_subscript0_share1_1 ; 
        x1x2x4x5x7_subscript0_share2_reg <= x1x2x4x5x7_subscript0_share2_1 ; 
        x1x3x4x6x7_subscript0_share1_reg <= x1x3x4x6x7_subscript0_share1_1 ; 
        x1x3x4x6x7_subscript0_share2_reg <= x1x3x4x6x7_subscript0_share2_1 ; 
        x1x3x5x6x7_subscript0_share1_reg <= x1x3x5x6x7_subscript0_share1_1 ; 
        x1x3x5x6x7_subscript0_share2_reg <= x1x3x5x6x7_subscript0_share2_1 ; 
        x1x4x5x6x7_subscript0_share1_reg <= x1x4x5x6x7_subscript0_share1_1 ; 
        x1x4x5x6x7_subscript0_share2_reg <= x1x4x5x6x7_subscript0_share2_1 ; 
        x2x3x5x6x7_subscript0_share1_reg <= x2x3x5x6x7_subscript0_share1_1 ; 
        x2x3x5x6x7_subscript0_share2_reg <= x2x3x5x6x7_subscript0_share2_1 ; 
        x3x4x5x6x7_subscript0_share1_reg <= x3x4x5x6x7_subscript0_share1_1 ; 
        x3x4x5x6x7_subscript0_share2_reg <= x3x4x5x6x7_subscript0_share2_1 ; 
        x0x1x2x5x6_subscript0_share1_reg <= x0x1x2x5x6_subscript0_share1_1 ; 
        x0x1x2x5x6_subscript0_share2_reg <= x0x1x2x5x6_subscript0_share2_1 ; 
        x0x1x3x4x5_subscript0_share1_reg <= x0x1x3x4x5_subscript0_share1_1 ; 
        x0x1x3x4x5_subscript0_share2_reg <= x0x1x3x4x5_subscript0_share2_1 ; 
        x0x1x4x5x7_subscript0_share1_reg <= x0x1x4x5x7_subscript0_share1_1 ; 
        x0x1x4x5x7_subscript0_share2_reg <= x0x1x4x5x7_subscript0_share2_1 ; 
        x0x2x3x5x6_subscript0_share1_reg <= x0x2x3x5x6_subscript0_share1_1 ; 
        x0x2x3x5x6_subscript0_share2_reg <= x0x2x3x5x6_subscript0_share2_1 ; 
        x1x2x3x4x7_subscript0_share1_reg <= x1x2x3x4x7_subscript0_share1_1 ; 
        x1x2x3x4x7_subscript0_share2_reg <= x1x2x3x4x7_subscript0_share2_1 ; 
        x0x1x2x3x4x6_subscript0_share1_reg <= x0x1x2x3x4x6_subscript0_share1_1 ; 
        x0x1x2x3x4x6_subscript0_share2_reg <= x0x1x2x3x4x6_subscript0_share2_1 ; 
        x0x1x2x3x4x7_subscript0_share1_reg <= x0x1x2x3x4x7_subscript0_share1_1 ; 
        x0x1x2x3x4x7_subscript0_share2_reg <= x0x1x2x3x4x7_subscript0_share2_1 ; 
        x0x1x2x3x5x7_subscript0_share1_reg <= x0x1x2x3x5x7_subscript0_share1_1 ; 
        x0x1x2x3x5x7_subscript0_share2_reg <= x0x1x2x3x5x7_subscript0_share2_1 ; 
        x0x1x2x3x6x7_subscript0_share1_reg <= x0x1x2x3x6x7_subscript0_share1_1 ; 
        x0x1x2x3x6x7_subscript0_share2_reg <= x0x1x2x3x6x7_subscript0_share2_1 ; 
        x0x1x2x4x5x7_subscript0_share1_reg <= x0x1x2x4x5x7_subscript0_share1_1 ; 
        x0x1x2x4x5x7_subscript0_share2_reg <= x0x1x2x4x5x7_subscript0_share2_1 ; 
        x0x1x2x5x6x7_subscript0_share1_reg <= x0x1x2x5x6x7_subscript0_share1_1 ; 
        x0x1x2x5x6x7_subscript0_share2_reg <= x0x1x2x5x6x7_subscript0_share2_1 ; 
        x0x1x3x4x6x7_subscript0_share1_reg <= x0x1x3x4x6x7_subscript0_share1_1 ; 
        x0x1x3x4x6x7_subscript0_share2_reg <= x0x1x3x4x6x7_subscript0_share2_1 ; 
        x0x1x4x5x6x7_subscript0_share1_reg <= x0x1x4x5x6x7_subscript0_share1_1 ; 
        x0x1x4x5x6x7_subscript0_share2_reg <= x0x1x4x5x6x7_subscript0_share2_1 ; 
        x0x2x3x4x5x6_subscript0_share1_reg <= x0x2x3x4x5x6_subscript0_share1_1 ; 
        x0x2x3x4x5x6_subscript0_share2_reg <= x0x2x3x4x5x6_subscript0_share2_1 ; 
        x0x2x3x4x5x7_subscript0_share1_reg <= x0x2x3x4x5x7_subscript0_share1_1 ; 
        x0x2x3x4x5x7_subscript0_share2_reg <= x0x2x3x4x5x7_subscript0_share2_1 ; 
        x0x2x3x5x6x7_subscript0_share1_reg <= x0x2x3x5x6x7_subscript0_share1_1 ; 
        x0x2x3x5x6x7_subscript0_share2_reg <= x0x2x3x5x6x7_subscript0_share2_1 ; 
        x1x2x3x4x6x7_subscript0_share1_reg <= x1x2x3x4x6x7_subscript0_share1_1 ; 
        x1x2x3x4x6x7_subscript0_share2_reg <= x1x2x3x4x6x7_subscript0_share2_1 ; 
        x1x2x4x5x6x7_subscript0_share1_reg <= x1x2x4x5x6x7_subscript0_share1_1 ; 
        x1x2x4x5x6x7_subscript0_share2_reg <= x1x2x4x5x6x7_subscript0_share2_1 ; 
        x1x3x4x5x6x7_subscript0_share1_reg <= x1x3x4x5x6x7_subscript0_share1_1 ; 
        x1x3x4x5x6x7_subscript0_share2_reg <= x1x3x4x5x6x7_subscript0_share2_1 ; 
        x2x3x4x5x6x7_subscript0_share1_reg <= x2x3x4x5x6x7_subscript0_share1_1 ; 
        x2x3x4x5x6x7_subscript0_share2_reg <= x2x3x4x5x6x7_subscript0_share2_1 ; 
        x0x1x2x3x5x6_subscript0_share1_reg <= x0x1x2x3x5x6_subscript0_share1_1 ; 
        x0x1x2x3x5x6_subscript0_share2_reg <= x0x1x2x3x5x6_subscript0_share2_1 ; 
        x0x1x2x4x6x7_subscript0_share1_reg <= x0x1x2x4x6x7_subscript0_share1_1 ; 
        x0x1x2x4x6x7_subscript0_share2_reg <= x0x1x2x4x6x7_subscript0_share2_1 ; 
        x0x1x3x4x5x6_subscript0_share1_reg <= x0x1x3x4x5x6_subscript0_share1_1 ; 
        x0x1x3x4x5x6_subscript0_share2_reg <= x0x1x3x4x5x6_subscript0_share2_1 ; 
        x0x2x3x4x6x7_subscript0_share1_reg <= x0x2x3x4x6x7_subscript0_share1_1 ; 
        x0x2x3x4x6x7_subscript0_share2_reg <= x0x2x3x4x6x7_subscript0_share2_1 ; 
        x1x2x3x4x5x6_subscript0_share1_reg <= x1x2x3x4x5x6_subscript0_share1_1 ; 
        x1x2x3x4x5x6_subscript0_share2_reg <= x1x2x3x4x5x6_subscript0_share2_1 ; 
        x1x2x3x5x6x7_subscript0_share1_reg <= x1x2x3x5x6x7_subscript0_share1_1 ; 
        x1x2x3x5x6x7_subscript0_share2_reg <= x1x2x3x5x6x7_subscript0_share2_1 ; 
        x0x1x2x3x4x5_subscript0_share1_reg <= x0x1x2x3x4x5_subscript0_share1_1 ; 
        x0x1x2x3x4x5_subscript0_share2_reg <= x0x1x2x3x4x5_subscript0_share2_1 ; 
        x0x1x2x4x5x6_subscript0_share1_reg <= x0x1x2x4x5x6_subscript0_share1_1 ; 
        x0x1x2x4x5x6_subscript0_share2_reg <= x0x1x2x4x5x6_subscript0_share2_1 ; 
        x0x1x3x4x5x7_subscript0_share1_reg <= x0x1x3x4x5x7_subscript0_share1_1 ; 
        x0x1x3x4x5x7_subscript0_share2_reg <= x0x1x3x4x5x7_subscript0_share2_1 ; 
        x0x1x3x5x6x7_subscript0_share1_reg <= x0x1x3x5x6x7_subscript0_share1_1 ; 
        x0x1x3x5x6x7_subscript0_share2_reg <= x0x1x3x5x6x7_subscript0_share2_1 ; 
        x0x2x4x5x6x7_subscript0_share1_reg <= x0x2x4x5x6x7_subscript0_share1_1 ; 
        x0x2x4x5x6x7_subscript0_share2_reg <= x0x2x4x5x6x7_subscript0_share2_1 ; 
        x1x2x3x4x5x7_subscript0_share1_reg <= x1x2x3x4x5x7_subscript0_share1_1 ; 
        x1x2x3x4x5x7_subscript0_share2_reg <= x1x2x3x4x5x7_subscript0_share2_1 ; 
        x0x3x4x5x6x7_subscript0_share1_reg <= x0x3x4x5x6x7_subscript0_share1_1 ; 
        x0x3x4x5x6x7_subscript0_share2_reg <= x0x3x4x5x6x7_subscript0_share2_1 ; 
        x0x1x2x3x4x6x7_subscript0_share1_reg <= x0x1x2x3x4x6x7_subscript0_share1_1 ; 
        x0x1x2x3x4x6x7_subscript0_share2_reg <= x0x1x2x3x4x6x7_subscript0_share2_1 ; 
        x0x1x2x4x5x6x7_subscript0_share1_reg <= x0x1x2x4x5x6x7_subscript0_share1_1 ; 
        x0x1x2x4x5x6x7_subscript0_share2_reg <= x0x1x2x4x5x6x7_subscript0_share2_1 ; 
        x0x2x3x4x5x6x7_subscript0_share1_reg <= x0x2x3x4x5x6x7_subscript0_share1_1 ; 
        x0x2x3x4x5x6x7_subscript0_share2_reg <= x0x2x3x4x5x6x7_subscript0_share2_1 ; 
        x0x1x2x3x5x6x7_subscript0_share1_reg <= x0x1x2x3x5x6x7_subscript0_share1_1 ; 
        x0x1x2x3x5x6x7_subscript0_share2_reg <= x0x1x2x3x5x6x7_subscript0_share2_1 ; 
        x0x1x3x4x5x6x7_subscript0_share1_reg <= x0x1x3x4x5x6x7_subscript0_share1_1 ; 
        x0x1x3x4x5x6x7_subscript0_share2_reg <= x0x1x3x4x5x6x7_subscript0_share2_1 ; 
        x1x2x3x4x5x6x7_subscript0_share1_reg <= x1x2x3x4x5x6x7_subscript0_share1_1 ; 
        x1x2x3x4x5x6x7_subscript0_share2_reg <= x1x2x3x4x5x6x7_subscript0_share2_1 ; 
        x0x1x2x3x4x5x6_subscript0_share1_reg <= x0x1x2x3x4x5x6_subscript0_share1_1 ; 
        x0x1x2x3x4x5x6_subscript0_share2_reg <= x0x1x2x3x4x5x6_subscript0_share2_1 ; 
        x0x1x2x3x4x5x7_subscript0_share1_reg <= x0x1x2x3x4x5x7_subscript0_share1_1 ; 
        x0x1x2x3x4x5x7_subscript0_share2_reg <= x0x1x2x3x4x5x7_subscript0_share2_1 ; 

end

wire [7:0] output_sbox_share1, output_sbox_share2, output_sbox;

assign output_sbox_share1 = { sbox_out1_share1, sbox_out2_share1, sbox_out3_share1, sbox_out4_share1, sbox_out5_share1, sbox_out6_share1, sbox_out7_share1, sbox_out8_share1};
assign output_sbox_share2 = { sbox_out1_share2, sbox_out2_share2, sbox_out3_share2, sbox_out4_share2, sbox_out5_share2, sbox_out6_share2, sbox_out7_share2, sbox_out8_share2};


assign sbox_output_share1 = output_sbox_share1; 
assign sbox_output_share2 = output_sbox_share2; 

endmodule
