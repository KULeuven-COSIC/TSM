`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:        COSIC, KU Leuven, Belgium
// Engineer:       Dilip Kumar S V
// Paper:          Higher-Order Time Sharing Masking
// Authors:        Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, 
//                 Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date:    02/22/2025
// Design Name:    Masked AES Round Function
// Module Name:    aes_round_function
// Description:    Implements the round function for AES with Time Sharing Masking. 
//                 This includes key addition, S-box transformation, row shifting, 
//                 column mixing, and the final output generation for both shares 
//                 of ciphertext.
// Dependencies:    AES S-box, two-dimensional array, XOR, and multiplexer modules.
// Revision:       0.01 - Initial version
//////////////////////////////////////////////////////////////////////////////////

module aes_round_function ( clk, reset, start,
rand_cycle1,rand_cycle2,
plaintext_share1, plaintext_share2, key_input_share1, key_input_share2, add_roundkey_share1, add_roundkey_share2,
out_done,ciphertext_share1,ciphertext_share2
);

input clk, reset,start;
input [608:1] rand_cycle1;
input [128:1] rand_cycle2;
input [128:1] plaintext_share1;
input [128:1] plaintext_share2;
input [128:1] key_input_share1;
input [128:1] key_input_share2;
input [128:1] add_roundkey_share1;
input [128:1] add_roundkey_share2;
output [128:1] ciphertext_share1;
output [128:1] ciphertext_share2;
output out_done;


wire [8:1] add_roundkey_share1_row1_col1, add_roundkey_share1_row1_col2, add_roundkey_share1_row1_col3, add_roundkey_share1_row1_col4, add_roundkey_share1_row2_col1, add_roundkey_share1_row2_col2, add_roundkey_share1_row2_col3, add_roundkey_share1_row2_col4, add_roundkey_share1_row3_col1, add_roundkey_share1_row3_col2, add_roundkey_share1_row3_col3, add_roundkey_share1_row3_col4, add_roundkey_share1_row4_col1, add_roundkey_share1_row4_col2, add_roundkey_share1_row4_col3, add_roundkey_share1_row4_col4 ;
wire [8:1] add_roundkey_share2_row1_col1, add_roundkey_share2_row1_col2, add_roundkey_share2_row1_col3, add_roundkey_share2_row1_col4, add_roundkey_share2_row2_col1, add_roundkey_share2_row2_col2, add_roundkey_share2_row2_col3, add_roundkey_share2_row2_col4, add_roundkey_share2_row3_col1, add_roundkey_share2_row3_col2, add_roundkey_share2_row3_col3, add_roundkey_share2_row3_col4, add_roundkey_share2_row4_col1, add_roundkey_share2_row4_col2, add_roundkey_share2_row4_col3, add_roundkey_share2_row4_col4 ;
wire [8:1] key_input_share1_row1_col1, key_input_share1_row1_col2, key_input_share1_row1_col3, key_input_share1_row1_col4, key_input_share1_row2_col1, key_input_share1_row2_col2, key_input_share1_row2_col3, key_input_share1_row2_col4, key_input_share1_row3_col1, key_input_share1_row3_col2, key_input_share1_row3_col3, key_input_share1_row3_col4, key_input_share1_row4_col1, key_input_share1_row4_col2, key_input_share1_row4_col3, key_input_share1_row4_col4 ;
wire [8:1] key_input_share2_row1_col1, key_input_share2_row1_col2, key_input_share2_row1_col3, key_input_share2_row1_col4, key_input_share2_row2_col1, key_input_share2_row2_col2, key_input_share2_row2_col3, key_input_share2_row2_col4, key_input_share2_row3_col1, key_input_share2_row3_col2, key_input_share2_row3_col3, key_input_share2_row3_col4, key_input_share2_row4_col1, key_input_share2_row4_col2, key_input_share2_row4_col3, key_input_share2_row4_col4 ;
wire [8:1] plaintext_share1_row1_col1, plaintext_share1_row1_col2, plaintext_share1_row1_col3, plaintext_share1_row1_col4, plaintext_share1_row2_col1, plaintext_share1_row2_col2, plaintext_share1_row2_col3, plaintext_share1_row2_col4, plaintext_share1_row3_col1, plaintext_share1_row3_col2, plaintext_share1_row3_col3, plaintext_share1_row3_col4, plaintext_share1_row4_col1, plaintext_share1_row4_col2, plaintext_share1_row4_col3, plaintext_share1_row4_col4 ;
wire [8:1] plaintext_share2_row1_col1, plaintext_share2_row1_col2, plaintext_share2_row1_col3, plaintext_share2_row1_col4, plaintext_share2_row2_col1, plaintext_share2_row2_col2, plaintext_share2_row2_col3, plaintext_share2_row2_col4, plaintext_share2_row3_col1, plaintext_share2_row3_col2, plaintext_share2_row3_col3, plaintext_share2_row3_col4, plaintext_share2_row4_col1, plaintext_share2_row4_col2, plaintext_share2_row4_col3, plaintext_share2_row4_col4 ;


two_dimension_array inst_two_dimension_array_rkey_share1(
add_roundkey_share1,
add_roundkey_share1_row1_col1, add_roundkey_share1_row1_col2, add_roundkey_share1_row1_col3, add_roundkey_share1_row1_col4, add_roundkey_share1_row2_col1, add_roundkey_share1_row2_col2, add_roundkey_share1_row2_col3, add_roundkey_share1_row2_col4, add_roundkey_share1_row3_col1, add_roundkey_share1_row3_col2, add_roundkey_share1_row3_col3, add_roundkey_share1_row3_col4, add_roundkey_share1_row4_col1, add_roundkey_share1_row4_col2, add_roundkey_share1_row4_col3, add_roundkey_share1_row4_col4 
);
two_dimension_array inst_two_dimension_array_rkey_share2(
add_roundkey_share2,
add_roundkey_share2_row1_col1, add_roundkey_share2_row1_col2, add_roundkey_share2_row1_col3, add_roundkey_share2_row1_col4, add_roundkey_share2_row2_col1, add_roundkey_share2_row2_col2, add_roundkey_share2_row2_col3, add_roundkey_share2_row2_col4, add_roundkey_share2_row3_col1, add_roundkey_share2_row3_col2, add_roundkey_share2_row3_col3, add_roundkey_share2_row3_col4, add_roundkey_share2_row4_col1, add_roundkey_share2_row4_col2, add_roundkey_share2_row4_col3, add_roundkey_share2_row4_col4 
);

two_dimension_array inst_two_dimension_array_inputkey_share1(
key_input_share1,
key_input_share1_row1_col1, key_input_share1_row1_col2, key_input_share1_row1_col3, key_input_share1_row1_col4, key_input_share1_row2_col1, key_input_share1_row2_col2, key_input_share1_row2_col3, key_input_share1_row2_col4, key_input_share1_row3_col1, key_input_share1_row3_col2, key_input_share1_row3_col3, key_input_share1_row3_col4, key_input_share1_row4_col1, key_input_share1_row4_col2, key_input_share1_row4_col3, key_input_share1_row4_col4 
);
two_dimension_array inst_two_dimension_array_inputkey_share2(
key_input_share2,
key_input_share2_row1_col1, key_input_share2_row1_col2, key_input_share2_row1_col3, key_input_share2_row1_col4, key_input_share2_row2_col1, key_input_share2_row2_col2, key_input_share2_row2_col3, key_input_share2_row2_col4, key_input_share2_row3_col1, key_input_share2_row3_col2, key_input_share2_row3_col3, key_input_share2_row3_col4, key_input_share2_row4_col1, key_input_share2_row4_col2, key_input_share2_row4_col3, key_input_share2_row4_col4 
);
two_dimension_array inst_two_dimension_array_plaintext_share1(
plaintext_share1,
plaintext_share1_row1_col1, plaintext_share1_row1_col2, plaintext_share1_row1_col3, plaintext_share1_row1_col4, plaintext_share1_row2_col1, plaintext_share1_row2_col2, plaintext_share1_row2_col3, plaintext_share1_row2_col4, plaintext_share1_row3_col1, plaintext_share1_row3_col2, plaintext_share1_row3_col3, plaintext_share1_row3_col4, plaintext_share1_row4_col1, plaintext_share1_row4_col2, plaintext_share1_row4_col3, plaintext_share1_row4_col4 
);
two_dimension_array inst_two_dimension_array_plaintext_share2(
plaintext_share2,
plaintext_share2_row1_col1, plaintext_share2_row1_col2, plaintext_share2_row1_col3, plaintext_share2_row1_col4, plaintext_share2_row2_col1, plaintext_share2_row2_col2, plaintext_share2_row2_col3, plaintext_share2_row2_col4, plaintext_share2_row3_col1, plaintext_share2_row3_col2, plaintext_share2_row3_col3, plaintext_share2_row3_col4, plaintext_share2_row4_col1, plaintext_share2_row4_col2, plaintext_share2_row4_col3, plaintext_share2_row4_col4 
);



// First round input 

wire [8:1] first_round_sbox_input_share1_row1_col1, first_round_sbox_input_share1_row1_col2, first_round_sbox_input_share1_row1_col3, first_round_sbox_input_share1_row1_col4, first_round_sbox_input_share1_row2_col1, first_round_sbox_input_share1_row2_col2, first_round_sbox_input_share1_row2_col3, first_round_sbox_input_share1_row2_col4, first_round_sbox_input_share1_row3_col1, first_round_sbox_input_share1_row3_col2, first_round_sbox_input_share1_row3_col3, first_round_sbox_input_share1_row3_col4, first_round_sbox_input_share1_row4_col1, first_round_sbox_input_share1_row4_col2, first_round_sbox_input_share1_row4_col3, first_round_sbox_input_share1_row4_col4 ;
wire [8:1] first_round_sbox_input_share2_row1_col1, first_round_sbox_input_share2_row1_col2, first_round_sbox_input_share2_row1_col3, first_round_sbox_input_share2_row1_col4, first_round_sbox_input_share2_row2_col1, first_round_sbox_input_share2_row2_col2, first_round_sbox_input_share2_row2_col3, first_round_sbox_input_share2_row2_col4, first_round_sbox_input_share2_row3_col1, first_round_sbox_input_share2_row3_col2, first_round_sbox_input_share2_row3_col3, first_round_sbox_input_share2_row3_col4, first_round_sbox_input_share2_row4_col1, first_round_sbox_input_share2_row4_col2, first_round_sbox_input_share2_row4_col3, first_round_sbox_input_share2_row4_col4 ;

two_dimension_xor inst_first_round_sbox_input_xor_share1 (
key_input_share1_row1_col1, key_input_share1_row1_col2, key_input_share1_row1_col3, key_input_share1_row1_col4, key_input_share1_row2_col1, key_input_share1_row2_col2, key_input_share1_row2_col3, key_input_share1_row2_col4, key_input_share1_row3_col1, key_input_share1_row3_col2, key_input_share1_row3_col3, key_input_share1_row3_col4, key_input_share1_row4_col1, key_input_share1_row4_col2, key_input_share1_row4_col3, key_input_share1_row4_col4 ,
plaintext_share1_row1_col1, plaintext_share1_row1_col2, plaintext_share1_row1_col3, plaintext_share1_row1_col4, plaintext_share1_row2_col1, plaintext_share1_row2_col2, plaintext_share1_row2_col3, plaintext_share1_row2_col4, plaintext_share1_row3_col1, plaintext_share1_row3_col2, plaintext_share1_row3_col3, plaintext_share1_row3_col4, plaintext_share1_row4_col1, plaintext_share1_row4_col2, plaintext_share1_row4_col3, plaintext_share1_row4_col4 ,
first_round_sbox_input_share1_row1_col1, first_round_sbox_input_share1_row1_col2, first_round_sbox_input_share1_row1_col3, first_round_sbox_input_share1_row1_col4, first_round_sbox_input_share1_row2_col1, first_round_sbox_input_share1_row2_col2, first_round_sbox_input_share1_row2_col3, first_round_sbox_input_share1_row2_col4, first_round_sbox_input_share1_row3_col1, first_round_sbox_input_share1_row3_col2, first_round_sbox_input_share1_row3_col3, first_round_sbox_input_share1_row3_col4, first_round_sbox_input_share1_row4_col1, first_round_sbox_input_share1_row4_col2, first_round_sbox_input_share1_row4_col3, first_round_sbox_input_share1_row4_col4 
);
two_dimension_xor inst_first_round_sbox_input_xor_share2 (
key_input_share2_row1_col1, key_input_share2_row1_col2, key_input_share2_row1_col3, key_input_share2_row1_col4, key_input_share2_row2_col1, key_input_share2_row2_col2, key_input_share2_row2_col3, key_input_share2_row2_col4, key_input_share2_row3_col1, key_input_share2_row3_col2, key_input_share2_row3_col3, key_input_share2_row3_col4, key_input_share2_row4_col1, key_input_share2_row4_col2, key_input_share2_row4_col3, key_input_share2_row4_col4 ,
plaintext_share2_row1_col1, plaintext_share2_row1_col2, plaintext_share2_row1_col3, plaintext_share2_row1_col4, plaintext_share2_row2_col1, plaintext_share2_row2_col2, plaintext_share2_row2_col3, plaintext_share2_row2_col4, plaintext_share2_row3_col1, plaintext_share2_row3_col2, plaintext_share2_row3_col3, plaintext_share2_row3_col4, plaintext_share2_row4_col1, plaintext_share2_row4_col2, plaintext_share2_row4_col3, plaintext_share2_row4_col4 ,
first_round_sbox_input_share2_row1_col1, first_round_sbox_input_share2_row1_col2, first_round_sbox_input_share2_row1_col3, first_round_sbox_input_share2_row1_col4, first_round_sbox_input_share2_row2_col1, first_round_sbox_input_share2_row2_col2, first_round_sbox_input_share2_row2_col3, first_round_sbox_input_share2_row2_col4, first_round_sbox_input_share2_row3_col1, first_round_sbox_input_share2_row3_col2, first_round_sbox_input_share2_row3_col3, first_round_sbox_input_share2_row3_col4, first_round_sbox_input_share2_row4_col1, first_round_sbox_input_share2_row4_col2, first_round_sbox_input_share2_row4_col3, first_round_sbox_input_share2_row4_col4 
);

wire [8:1] sbox_input_share1_row1_col1, sbox_input_share1_row1_col2, sbox_input_share1_row1_col3, sbox_input_share1_row1_col4, sbox_input_share1_row2_col1, sbox_input_share1_row2_col2, sbox_input_share1_row2_col3, sbox_input_share1_row2_col4, sbox_input_share1_row3_col1, sbox_input_share1_row3_col2, sbox_input_share1_row3_col3, sbox_input_share1_row3_col4, sbox_input_share1_row4_col1, sbox_input_share1_row4_col2, sbox_input_share1_row4_col3, sbox_input_share1_row4_col4 ;
wire [8:1] sbox_input_share2_row1_col1, sbox_input_share2_row1_col2, sbox_input_share2_row1_col3, sbox_input_share2_row1_col4, sbox_input_share2_row2_col1, sbox_input_share2_row2_col2, sbox_input_share2_row2_col3, sbox_input_share2_row2_col4, sbox_input_share2_row3_col1, sbox_input_share2_row3_col2, sbox_input_share2_row3_col3, sbox_input_share2_row3_col4, sbox_input_share2_row4_col1, sbox_input_share2_row4_col2, sbox_input_share2_row4_col3, sbox_input_share2_row4_col4 ;
wire [8:1] next_state_share1_row1_col1, next_state_share1_row1_col2, next_state_share1_row1_col3, next_state_share1_row1_col4, next_state_share1_row2_col1, next_state_share1_row2_col2, next_state_share1_row2_col3, next_state_share1_row2_col4, next_state_share1_row3_col1, next_state_share1_row3_col2, next_state_share1_row3_col3, next_state_share1_row3_col4, next_state_share1_row4_col1, next_state_share1_row4_col2, next_state_share1_row4_col3, next_state_share1_row4_col4 ;
wire [8:1] next_state_share2_row1_col1, next_state_share2_row1_col2, next_state_share2_row1_col3, next_state_share2_row1_col4, next_state_share2_row2_col1, next_state_share2_row2_col2, next_state_share2_row2_col3, next_state_share2_row2_col4, next_state_share2_row3_col1, next_state_share2_row3_col2, next_state_share2_row3_col3, next_state_share2_row3_col4, next_state_share2_row4_col1, next_state_share2_row4_col2, next_state_share2_row4_col3, next_state_share2_row4_col4 ;

reg select_first_round, select_final_round;

wire [8:1] mixed_sbox_output_share1_row1_col1, mixed_sbox_output_share1_row1_col2, mixed_sbox_output_share1_row1_col3, mixed_sbox_output_share1_row1_col4, mixed_sbox_output_share1_row2_col1, mixed_sbox_output_share1_row2_col2, mixed_sbox_output_share1_row2_col3, mixed_sbox_output_share1_row2_col4, mixed_sbox_output_share1_row3_col1, mixed_sbox_output_share1_row3_col2, mixed_sbox_output_share1_row3_col3, mixed_sbox_output_share1_row3_col4, mixed_sbox_output_share1_row4_col1, mixed_sbox_output_share1_row4_col2, mixed_sbox_output_share1_row4_col3, mixed_sbox_output_share1_row4_col4 ;
wire [8:1] mixed_sbox_output_share2_row1_col1, mixed_sbox_output_share2_row1_col2, mixed_sbox_output_share2_row1_col3, mixed_sbox_output_share2_row1_col4, mixed_sbox_output_share2_row2_col1, mixed_sbox_output_share2_row2_col2, mixed_sbox_output_share2_row2_col3, mixed_sbox_output_share2_row2_col4, mixed_sbox_output_share2_row3_col1, mixed_sbox_output_share2_row3_col2, mixed_sbox_output_share2_row3_col3, mixed_sbox_output_share2_row3_col4, mixed_sbox_output_share2_row4_col1, mixed_sbox_output_share2_row4_col2, mixed_sbox_output_share2_row4_col3, mixed_sbox_output_share2_row4_col4 ;

two_dimension_mux inst_state_reg_share1_mux(
select_first_round, 
first_round_sbox_input_share1_row1_col1, first_round_sbox_input_share1_row1_col2, first_round_sbox_input_share1_row1_col3, first_round_sbox_input_share1_row1_col4, first_round_sbox_input_share1_row2_col1, first_round_sbox_input_share1_row2_col2, first_round_sbox_input_share1_row2_col3, first_round_sbox_input_share1_row2_col4, first_round_sbox_input_share1_row3_col1, first_round_sbox_input_share1_row3_col2, first_round_sbox_input_share1_row3_col3, first_round_sbox_input_share1_row3_col4, first_round_sbox_input_share1_row4_col1, first_round_sbox_input_share1_row4_col2, first_round_sbox_input_share1_row4_col3, first_round_sbox_input_share1_row4_col4 ,
next_state_share1_row1_col1, next_state_share1_row1_col2, next_state_share1_row1_col3, next_state_share1_row1_col4, next_state_share1_row2_col1, next_state_share1_row2_col2, next_state_share1_row2_col3, next_state_share1_row2_col4, next_state_share1_row3_col1, next_state_share1_row3_col2, next_state_share1_row3_col3, next_state_share1_row3_col4, next_state_share1_row4_col1, next_state_share1_row4_col2, next_state_share1_row4_col3, next_state_share1_row4_col4 ,
sbox_input_share1_row1_col1, sbox_input_share1_row1_col2, sbox_input_share1_row1_col3, sbox_input_share1_row1_col4, sbox_input_share1_row2_col1, sbox_input_share1_row2_col2, sbox_input_share1_row2_col3, sbox_input_share1_row2_col4, sbox_input_share1_row3_col1, sbox_input_share1_row3_col2, sbox_input_share1_row3_col3, sbox_input_share1_row3_col4, sbox_input_share1_row4_col1, sbox_input_share1_row4_col2, sbox_input_share1_row4_col3, sbox_input_share1_row4_col4 
);
two_dimension_mux inst_state_reg_share2_mux(
select_first_round, 
first_round_sbox_input_share2_row1_col1, first_round_sbox_input_share2_row1_col2, first_round_sbox_input_share2_row1_col3, first_round_sbox_input_share2_row1_col4, first_round_sbox_input_share2_row2_col1, first_round_sbox_input_share2_row2_col2, first_round_sbox_input_share2_row2_col3, first_round_sbox_input_share2_row2_col4, first_round_sbox_input_share2_row3_col1, first_round_sbox_input_share2_row3_col2, first_round_sbox_input_share2_row3_col3, first_round_sbox_input_share2_row3_col4, first_round_sbox_input_share2_row4_col1, first_round_sbox_input_share2_row4_col2, first_round_sbox_input_share2_row4_col3, first_round_sbox_input_share2_row4_col4 ,
next_state_share2_row1_col1, next_state_share2_row1_col2, next_state_share2_row1_col3, next_state_share2_row1_col4, next_state_share2_row2_col1, next_state_share2_row2_col2, next_state_share2_row2_col3, next_state_share2_row2_col4, next_state_share2_row3_col1, next_state_share2_row3_col2, next_state_share2_row3_col3, next_state_share2_row3_col4, next_state_share2_row4_col1, next_state_share2_row4_col2, next_state_share2_row4_col3, next_state_share2_row4_col4 ,
sbox_input_share2_row1_col1, sbox_input_share2_row1_col2, sbox_input_share2_row1_col3, sbox_input_share2_row1_col4, sbox_input_share2_row2_col1, sbox_input_share2_row2_col2, sbox_input_share2_row2_col3, sbox_input_share2_row2_col4, sbox_input_share2_row3_col1, sbox_input_share2_row3_col2, sbox_input_share2_row3_col3, sbox_input_share2_row3_col4, sbox_input_share2_row4_col1, sbox_input_share2_row4_col2, sbox_input_share2_row4_col3, sbox_input_share2_row4_col4 
);



wire [38:1] rand_cycle1_row1_col1 ,rand_cycle1_row1_col2 ,rand_cycle1_row1_col3 ,rand_cycle1_row1_col4 ,rand_cycle1_row2_col1 ,rand_cycle1_row2_col2 ,rand_cycle1_row2_col3 ,rand_cycle1_row2_col4 ,rand_cycle1_row3_col1 ,rand_cycle1_row3_col2 ,rand_cycle1_row3_col3 ,rand_cycle1_row3_col4 ,rand_cycle1_row4_col1 ,rand_cycle1_row4_col2 ,rand_cycle1_row4_col3 ,rand_cycle1_row4_col4 ;
wire [8:1]  rand_cycle2_row1_col1 ,rand_cycle2_row1_col2 ,rand_cycle2_row1_col3 ,rand_cycle2_row1_col4 ,rand_cycle2_row2_col1 ,rand_cycle2_row2_col2 ,rand_cycle2_row2_col3 ,rand_cycle2_row2_col4 ,rand_cycle2_row3_col1 ,rand_cycle2_row3_col2 ,rand_cycle2_row3_col3 ,rand_cycle2_row3_col4 ,rand_cycle2_row4_col1 ,rand_cycle2_row4_col2 ,rand_cycle2_row4_col3 ,rand_cycle2_row4_col4 ;
wire [8:1]  sbox_output_share1_row1_col1 ,sbox_output_share1_row1_col2 ,sbox_output_share1_row1_col3 ,sbox_output_share1_row1_col4 ,sbox_output_share1_row2_col1 ,sbox_output_share1_row2_col2 ,sbox_output_share1_row2_col3 ,sbox_output_share1_row2_col4 ,sbox_output_share1_row3_col1 ,sbox_output_share1_row3_col2 ,sbox_output_share1_row3_col3 ,sbox_output_share1_row3_col4 ,sbox_output_share1_row4_col1 ,sbox_output_share1_row4_col2 ,sbox_output_share1_row4_col3 ,sbox_output_share1_row4_col4 ;
wire [8:1]  sbox_output_share2_row1_col1 ,sbox_output_share2_row1_col2 ,sbox_output_share2_row1_col3 ,sbox_output_share2_row1_col4 ,sbox_output_share2_row2_col1 ,sbox_output_share2_row2_col2 ,sbox_output_share2_row2_col3 ,sbox_output_share2_row2_col4 ,sbox_output_share2_row3_col1 ,sbox_output_share2_row3_col2 ,sbox_output_share2_row3_col3 ,sbox_output_share2_row3_col4 ,sbox_output_share2_row4_col1 ,sbox_output_share2_row4_col2 ,sbox_output_share2_row4_col3 ,sbox_output_share2_row4_col4 ;

assign rand_cycle1_row1_col1 = rand_cycle1[38:1]    ;
assign rand_cycle1_row1_col2 = rand_cycle1[76:39]    ;
assign rand_cycle1_row1_col3 = rand_cycle1[114:77]    ;
assign rand_cycle1_row1_col4 = rand_cycle1[152:115]    ;
assign rand_cycle1_row2_col1 = rand_cycle1[190:153]    ;
assign rand_cycle1_row2_col2 = rand_cycle1[228:191]    ;
assign rand_cycle1_row2_col3 = rand_cycle1[266:229]    ;
assign rand_cycle1_row2_col4 = rand_cycle1[304:267]    ;
assign rand_cycle1_row3_col1 = rand_cycle1[342:305]    ;
assign rand_cycle1_row3_col2 = rand_cycle1[380:343]    ;
assign rand_cycle1_row3_col3 = rand_cycle1[418:381]    ;
assign rand_cycle1_row3_col4 = rand_cycle1[456:419]    ;
assign rand_cycle1_row4_col1 = rand_cycle1[494:457]    ;
assign rand_cycle1_row4_col2 = rand_cycle1[532:495]    ;
assign rand_cycle1_row4_col3 = rand_cycle1[570:533]    ;
assign rand_cycle1_row4_col4 = rand_cycle1[608:571]    ;

assign rand_cycle2_row1_col1 = rand_cycle2[8:1]    ;
assign rand_cycle2_row1_col2 = rand_cycle2[16:9]    ;
assign rand_cycle2_row1_col3 = rand_cycle2[24:17]    ;
assign rand_cycle2_row1_col4 = rand_cycle2[32:25]    ;
assign rand_cycle2_row2_col1 = rand_cycle2[40:33]    ;
assign rand_cycle2_row2_col2 = rand_cycle2[48:41]    ;
assign rand_cycle2_row2_col3 = rand_cycle2[56:49]    ;
assign rand_cycle2_row2_col4 = rand_cycle2[64:57]    ;
assign rand_cycle2_row3_col1 = rand_cycle2[72:65]    ;
assign rand_cycle2_row3_col2 = rand_cycle2[80:73]    ;
assign rand_cycle2_row3_col3 = rand_cycle2[88:81]    ;
assign rand_cycle2_row3_col4 = rand_cycle2[96:89]    ;
assign rand_cycle2_row4_col1 = rand_cycle2[104:97]    ;
assign rand_cycle2_row4_col2 = rand_cycle2[112:105]    ;
assign rand_cycle2_row4_col3 = rand_cycle2[120:113]    ;
assign rand_cycle2_row4_col4 = rand_cycle2[128:121]    ;


reg enable_sbox_cycle1, enable_sbox_cycle2 ;


AES_sbox_twocycle_firstorder inst_sbox_row1_col1 ( clk, rand_cycle1_row1_col1, rand_cycle2_row1_col1,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row1_col1,  sbox_input_share2_row1_col1,    sbox_output_share1_row1_col1,  sbox_output_share2_row1_col1 );
AES_sbox_twocycle_firstorder inst_sbox_row2_col1 ( clk, rand_cycle1_row2_col1, rand_cycle2_row2_col1,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row2_col1,  sbox_input_share2_row2_col1,    sbox_output_share1_row2_col1,  sbox_output_share2_row2_col1 );
AES_sbox_twocycle_firstorder inst_sbox_row3_col1 ( clk, rand_cycle1_row3_col1, rand_cycle2_row3_col1,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row3_col1,  sbox_input_share2_row3_col1,    sbox_output_share1_row3_col1,  sbox_output_share2_row3_col1 );
AES_sbox_twocycle_firstorder inst_sbox_row4_col1 ( clk, rand_cycle1_row4_col1, rand_cycle2_row4_col1,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row4_col1,  sbox_input_share2_row4_col1,    sbox_output_share1_row4_col1,  sbox_output_share2_row4_col1 );
AES_sbox_twocycle_firstorder inst_sbox_row1_col2 ( clk, rand_cycle1_row1_col2, rand_cycle2_row1_col2,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row1_col2,  sbox_input_share2_row1_col2,    sbox_output_share1_row1_col2,  sbox_output_share2_row1_col2 );
AES_sbox_twocycle_firstorder inst_sbox_row2_col2 ( clk, rand_cycle1_row2_col2, rand_cycle2_row2_col2,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row2_col2,  sbox_input_share2_row2_col2,    sbox_output_share1_row2_col2,  sbox_output_share2_row2_col2 );
AES_sbox_twocycle_firstorder inst_sbox_row3_col2 ( clk, rand_cycle1_row3_col2, rand_cycle2_row3_col2,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row3_col2,  sbox_input_share2_row3_col2,    sbox_output_share1_row3_col2,  sbox_output_share2_row3_col2 );
AES_sbox_twocycle_firstorder inst_sbox_row4_col2 ( clk, rand_cycle1_row4_col2, rand_cycle2_row4_col2,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row4_col2,  sbox_input_share2_row4_col2,    sbox_output_share1_row4_col2,  sbox_output_share2_row4_col2 );
AES_sbox_twocycle_firstorder inst_sbox_row1_col3 ( clk, rand_cycle1_row1_col3, rand_cycle2_row1_col3,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row1_col3,  sbox_input_share2_row1_col3,    sbox_output_share1_row1_col3,  sbox_output_share2_row1_col3 );
AES_sbox_twocycle_firstorder inst_sbox_row2_col3 ( clk, rand_cycle1_row2_col3, rand_cycle2_row2_col3,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row2_col3,  sbox_input_share2_row2_col3,    sbox_output_share1_row2_col3,  sbox_output_share2_row2_col3 );
AES_sbox_twocycle_firstorder inst_sbox_row3_col3 ( clk, rand_cycle1_row3_col3, rand_cycle2_row3_col3,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row3_col3,  sbox_input_share2_row3_col3,    sbox_output_share1_row3_col3,  sbox_output_share2_row3_col3 );
AES_sbox_twocycle_firstorder inst_sbox_row4_col3 ( clk, rand_cycle1_row4_col3, rand_cycle2_row4_col3,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row4_col3,  sbox_input_share2_row4_col3,    sbox_output_share1_row4_col3,  sbox_output_share2_row4_col3 );
AES_sbox_twocycle_firstorder inst_sbox_row1_col4 ( clk, rand_cycle1_row1_col4, rand_cycle2_row1_col4,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row1_col4,  sbox_input_share2_row1_col4,    sbox_output_share1_row1_col4,  sbox_output_share2_row1_col4 );
AES_sbox_twocycle_firstorder inst_sbox_row2_col4 ( clk, rand_cycle1_row2_col4, rand_cycle2_row2_col4,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row2_col4,  sbox_input_share2_row2_col4,    sbox_output_share1_row2_col4,  sbox_output_share2_row2_col4 );
AES_sbox_twocycle_firstorder inst_sbox_row3_col4 ( clk, rand_cycle1_row3_col4, rand_cycle2_row3_col4,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row3_col4,  sbox_input_share2_row3_col4,    sbox_output_share1_row3_col4,  sbox_output_share2_row3_col4 );
AES_sbox_twocycle_firstorder inst_sbox_row4_col4 ( clk, rand_cycle1_row4_col4, rand_cycle2_row4_col4,	reset, enable_sbox_cycle1,	reset, enable_sbox_cycle2,	sbox_input_share1_row4_col4,  sbox_input_share2_row4_col4,    sbox_output_share1_row4_col4,  sbox_output_share2_row4_col4 );


wire [8:1] shifted_sbox_output_share1_row1_col1, shifted_sbox_output_share1_row1_col2, shifted_sbox_output_share1_row1_col3, shifted_sbox_output_share1_row1_col4, shifted_sbox_output_share1_row2_col1, shifted_sbox_output_share1_row2_col2, shifted_sbox_output_share1_row2_col3, shifted_sbox_output_share1_row2_col4, shifted_sbox_output_share1_row3_col1, shifted_sbox_output_share1_row3_col2, shifted_sbox_output_share1_row3_col3, shifted_sbox_output_share1_row3_col4, shifted_sbox_output_share1_row4_col1, shifted_sbox_output_share1_row4_col2, shifted_sbox_output_share1_row4_col3, shifted_sbox_output_share1_row4_col4 ;
wire [8:1] shifted_sbox_output_share2_row1_col1, shifted_sbox_output_share2_row1_col2, shifted_sbox_output_share2_row1_col3, shifted_sbox_output_share2_row1_col4, shifted_sbox_output_share2_row2_col1, shifted_sbox_output_share2_row2_col2, shifted_sbox_output_share2_row2_col3, shifted_sbox_output_share2_row2_col4, shifted_sbox_output_share2_row3_col1, shifted_sbox_output_share2_row3_col2, shifted_sbox_output_share2_row3_col3, shifted_sbox_output_share2_row3_col4, shifted_sbox_output_share2_row4_col1, shifted_sbox_output_share2_row4_col2, shifted_sbox_output_share2_row4_col3, shifted_sbox_output_share2_row4_col4 ;

aes_shift_row inst_shift_row_share1 (
sbox_output_share1_row1_col1, sbox_output_share1_row1_col2, sbox_output_share1_row1_col3, sbox_output_share1_row1_col4, sbox_output_share1_row2_col1, sbox_output_share1_row2_col2, sbox_output_share1_row2_col3, sbox_output_share1_row2_col4, sbox_output_share1_row3_col1, sbox_output_share1_row3_col2, sbox_output_share1_row3_col3, sbox_output_share1_row3_col4, sbox_output_share1_row4_col1, sbox_output_share1_row4_col2, sbox_output_share1_row4_col3, sbox_output_share1_row4_col4 ,
shifted_sbox_output_share1_row1_col1, shifted_sbox_output_share1_row1_col2, shifted_sbox_output_share1_row1_col3, shifted_sbox_output_share1_row1_col4, shifted_sbox_output_share1_row2_col1, shifted_sbox_output_share1_row2_col2, shifted_sbox_output_share1_row2_col3, shifted_sbox_output_share1_row2_col4, shifted_sbox_output_share1_row3_col1, shifted_sbox_output_share1_row3_col2, shifted_sbox_output_share1_row3_col3, shifted_sbox_output_share1_row3_col4, shifted_sbox_output_share1_row4_col1, shifted_sbox_output_share1_row4_col2, shifted_sbox_output_share1_row4_col3, shifted_sbox_output_share1_row4_col4 
);
aes_shift_row inst_shift_row_share2 (
sbox_output_share2_row1_col1, sbox_output_share2_row1_col2, sbox_output_share2_row1_col3, sbox_output_share2_row1_col4, sbox_output_share2_row2_col1, sbox_output_share2_row2_col2, sbox_output_share2_row2_col3, sbox_output_share2_row2_col4, sbox_output_share2_row3_col1, sbox_output_share2_row3_col2, sbox_output_share2_row3_col3, sbox_output_share2_row3_col4, sbox_output_share2_row4_col1, sbox_output_share2_row4_col2, sbox_output_share2_row4_col3, sbox_output_share2_row4_col4 ,
shifted_sbox_output_share2_row1_col1, shifted_sbox_output_share2_row1_col2, shifted_sbox_output_share2_row1_col3, shifted_sbox_output_share2_row1_col4, shifted_sbox_output_share2_row2_col1, shifted_sbox_output_share2_row2_col2, shifted_sbox_output_share2_row2_col3, shifted_sbox_output_share2_row2_col4, shifted_sbox_output_share2_row3_col1, shifted_sbox_output_share2_row3_col2, shifted_sbox_output_share2_row3_col3, shifted_sbox_output_share2_row3_col4, shifted_sbox_output_share2_row4_col1, shifted_sbox_output_share2_row4_col2, shifted_sbox_output_share2_row4_col3, shifted_sbox_output_share2_row4_col4 
);

aes_mixcolumn inst_col1_mixcolumn_share1 (shifted_sbox_output_share1_row1_col1,shifted_sbox_output_share1_row2_col1,shifted_sbox_output_share1_row3_col1,shifted_sbox_output_share1_row4_col1 , mixed_sbox_output_share1_row1_col1,mixed_sbox_output_share1_row2_col1,mixed_sbox_output_share1_row3_col1,mixed_sbox_output_share1_row4_col1 );
aes_mixcolumn inst_col2_mixcolumn_share1 (shifted_sbox_output_share1_row1_col2,shifted_sbox_output_share1_row2_col2,shifted_sbox_output_share1_row3_col2,shifted_sbox_output_share1_row4_col2 , mixed_sbox_output_share1_row1_col2,mixed_sbox_output_share1_row2_col2,mixed_sbox_output_share1_row3_col2,mixed_sbox_output_share1_row4_col2 );
aes_mixcolumn inst_col3_mixcolumn_share1 (shifted_sbox_output_share1_row1_col3,shifted_sbox_output_share1_row2_col3,shifted_sbox_output_share1_row3_col3,shifted_sbox_output_share1_row4_col3 , mixed_sbox_output_share1_row1_col3,mixed_sbox_output_share1_row2_col3,mixed_sbox_output_share1_row3_col3,mixed_sbox_output_share1_row4_col3 );
aes_mixcolumn inst_col4_mixcolumn_share1 (shifted_sbox_output_share1_row1_col4,shifted_sbox_output_share1_row2_col4,shifted_sbox_output_share1_row3_col4,shifted_sbox_output_share1_row4_col4 , mixed_sbox_output_share1_row1_col4,mixed_sbox_output_share1_row2_col4,mixed_sbox_output_share1_row3_col4,mixed_sbox_output_share1_row4_col4 );
aes_mixcolumn inst_col1_mixcolumn_share2 (shifted_sbox_output_share2_row1_col1,shifted_sbox_output_share2_row2_col1,shifted_sbox_output_share2_row3_col1,shifted_sbox_output_share2_row4_col1 , mixed_sbox_output_share2_row1_col1,mixed_sbox_output_share2_row2_col1,mixed_sbox_output_share2_row3_col1,mixed_sbox_output_share2_row4_col1 );
aes_mixcolumn inst_col2_mixcolumn_share2 (shifted_sbox_output_share2_row1_col2,shifted_sbox_output_share2_row2_col2,shifted_sbox_output_share2_row3_col2,shifted_sbox_output_share2_row4_col2 , mixed_sbox_output_share2_row1_col2,mixed_sbox_output_share2_row2_col2,mixed_sbox_output_share2_row3_col2,mixed_sbox_output_share2_row4_col2 );
aes_mixcolumn inst_col3_mixcolumn_share2 (shifted_sbox_output_share2_row1_col3,shifted_sbox_output_share2_row2_col3,shifted_sbox_output_share2_row3_col3,shifted_sbox_output_share2_row4_col3 , mixed_sbox_output_share2_row1_col3,mixed_sbox_output_share2_row2_col3,mixed_sbox_output_share2_row3_col3,mixed_sbox_output_share2_row4_col3 );
aes_mixcolumn inst_col4_mixcolumn_share2 (shifted_sbox_output_share2_row1_col4,shifted_sbox_output_share2_row2_col4,shifted_sbox_output_share2_row3_col4,shifted_sbox_output_share2_row4_col4 , mixed_sbox_output_share2_row1_col4,mixed_sbox_output_share2_row2_col4,mixed_sbox_output_share2_row3_col4,mixed_sbox_output_share2_row4_col4 );

wire [8:1] final_sbox_output_share1_row1_col1, final_sbox_output_share1_row1_col2, final_sbox_output_share1_row1_col3, final_sbox_output_share1_row1_col4, final_sbox_output_share1_row2_col1, final_sbox_output_share1_row2_col2, final_sbox_output_share1_row2_col3, final_sbox_output_share1_row2_col4, final_sbox_output_share1_row3_col1, final_sbox_output_share1_row3_col2, final_sbox_output_share1_row3_col3, final_sbox_output_share1_row3_col4, final_sbox_output_share1_row4_col1, final_sbox_output_share1_row4_col2, final_sbox_output_share1_row4_col3, final_sbox_output_share1_row4_col4 ;
wire [8:1] final_sbox_output_share2_row1_col1, final_sbox_output_share2_row1_col2, final_sbox_output_share2_row1_col3, final_sbox_output_share2_row1_col4, final_sbox_output_share2_row2_col1, final_sbox_output_share2_row2_col2, final_sbox_output_share2_row2_col3, final_sbox_output_share2_row2_col4, final_sbox_output_share2_row3_col1, final_sbox_output_share2_row3_col2, final_sbox_output_share2_row3_col3, final_sbox_output_share2_row3_col4, final_sbox_output_share2_row4_col1, final_sbox_output_share2_row4_col2, final_sbox_output_share2_row4_col3, final_sbox_output_share2_row4_col4 ;

two_dimension_mux inst_final_round_share1_mux(
select_final_round, 
shifted_sbox_output_share1_row1_col1, shifted_sbox_output_share1_row1_col2, shifted_sbox_output_share1_row1_col3, shifted_sbox_output_share1_row1_col4, shifted_sbox_output_share1_row2_col1, shifted_sbox_output_share1_row2_col2, shifted_sbox_output_share1_row2_col3, shifted_sbox_output_share1_row2_col4, shifted_sbox_output_share1_row3_col1, shifted_sbox_output_share1_row3_col2, shifted_sbox_output_share1_row3_col3, shifted_sbox_output_share1_row3_col4, shifted_sbox_output_share1_row4_col1, shifted_sbox_output_share1_row4_col2, shifted_sbox_output_share1_row4_col3, shifted_sbox_output_share1_row4_col4 ,
mixed_sbox_output_share1_row1_col1, mixed_sbox_output_share1_row1_col2, mixed_sbox_output_share1_row1_col3, mixed_sbox_output_share1_row1_col4, mixed_sbox_output_share1_row2_col1, mixed_sbox_output_share1_row2_col2, mixed_sbox_output_share1_row2_col3, mixed_sbox_output_share1_row2_col4, mixed_sbox_output_share1_row3_col1, mixed_sbox_output_share1_row3_col2, mixed_sbox_output_share1_row3_col3, mixed_sbox_output_share1_row3_col4, mixed_sbox_output_share1_row4_col1, mixed_sbox_output_share1_row4_col2, mixed_sbox_output_share1_row4_col3, mixed_sbox_output_share1_row4_col4 ,
final_sbox_output_share1_row1_col1, final_sbox_output_share1_row1_col2, final_sbox_output_share1_row1_col3, final_sbox_output_share1_row1_col4, final_sbox_output_share1_row2_col1, final_sbox_output_share1_row2_col2, final_sbox_output_share1_row2_col3, final_sbox_output_share1_row2_col4, final_sbox_output_share1_row3_col1, final_sbox_output_share1_row3_col2, final_sbox_output_share1_row3_col3, final_sbox_output_share1_row3_col4, final_sbox_output_share1_row4_col1, final_sbox_output_share1_row4_col2, final_sbox_output_share1_row4_col3, final_sbox_output_share1_row4_col4 
);
two_dimension_mux inst_final_round_share2_mux(
select_final_round, 
shifted_sbox_output_share2_row1_col1, shifted_sbox_output_share2_row1_col2, shifted_sbox_output_share2_row1_col3, shifted_sbox_output_share2_row1_col4, shifted_sbox_output_share2_row2_col1, shifted_sbox_output_share2_row2_col2, shifted_sbox_output_share2_row2_col3, shifted_sbox_output_share2_row2_col4, shifted_sbox_output_share2_row3_col1, shifted_sbox_output_share2_row3_col2, shifted_sbox_output_share2_row3_col3, shifted_sbox_output_share2_row3_col4, shifted_sbox_output_share2_row4_col1, shifted_sbox_output_share2_row4_col2, shifted_sbox_output_share2_row4_col3, shifted_sbox_output_share2_row4_col4 ,
mixed_sbox_output_share2_row1_col1, mixed_sbox_output_share2_row1_col2, mixed_sbox_output_share2_row1_col3, mixed_sbox_output_share2_row1_col4, mixed_sbox_output_share2_row2_col1, mixed_sbox_output_share2_row2_col2, mixed_sbox_output_share2_row2_col3, mixed_sbox_output_share2_row2_col4, mixed_sbox_output_share2_row3_col1, mixed_sbox_output_share2_row3_col2, mixed_sbox_output_share2_row3_col3, mixed_sbox_output_share2_row3_col4, mixed_sbox_output_share2_row4_col1, mixed_sbox_output_share2_row4_col2, mixed_sbox_output_share2_row4_col3, mixed_sbox_output_share2_row4_col4 ,
final_sbox_output_share2_row1_col1, final_sbox_output_share2_row1_col2, final_sbox_output_share2_row1_col3, final_sbox_output_share2_row1_col4, final_sbox_output_share2_row2_col1, final_sbox_output_share2_row2_col2, final_sbox_output_share2_row2_col3, final_sbox_output_share2_row2_col4, final_sbox_output_share2_row3_col1, final_sbox_output_share2_row3_col2, final_sbox_output_share2_row3_col3, final_sbox_output_share2_row3_col4, final_sbox_output_share2_row4_col1, final_sbox_output_share2_row4_col2, final_sbox_output_share2_row4_col3, final_sbox_output_share2_row4_col4 
);

two_dimension_xor inst_next_round_sbox_input_xor_share1 (
add_roundkey_share1_row1_col1, add_roundkey_share1_row1_col2, add_roundkey_share1_row1_col3, add_roundkey_share1_row1_col4, add_roundkey_share1_row2_col1, add_roundkey_share1_row2_col2, add_roundkey_share1_row2_col3, add_roundkey_share1_row2_col4, add_roundkey_share1_row3_col1, add_roundkey_share1_row3_col2, add_roundkey_share1_row3_col3, add_roundkey_share1_row3_col4, add_roundkey_share1_row4_col1, add_roundkey_share1_row4_col2, add_roundkey_share1_row4_col3, add_roundkey_share1_row4_col4 ,
final_sbox_output_share1_row1_col1, final_sbox_output_share1_row1_col2, final_sbox_output_share1_row1_col3, final_sbox_output_share1_row1_col4, final_sbox_output_share1_row2_col1, final_sbox_output_share1_row2_col2, final_sbox_output_share1_row2_col3, final_sbox_output_share1_row2_col4, final_sbox_output_share1_row3_col1, final_sbox_output_share1_row3_col2, final_sbox_output_share1_row3_col3, final_sbox_output_share1_row3_col4, final_sbox_output_share1_row4_col1, final_sbox_output_share1_row4_col2, final_sbox_output_share1_row4_col3, final_sbox_output_share1_row4_col4 ,
next_state_share1_row1_col1, next_state_share1_row1_col2, next_state_share1_row1_col3, next_state_share1_row1_col4, next_state_share1_row2_col1, next_state_share1_row2_col2, next_state_share1_row2_col3, next_state_share1_row2_col4, next_state_share1_row3_col1, next_state_share1_row3_col2, next_state_share1_row3_col3, next_state_share1_row3_col4, next_state_share1_row4_col1, next_state_share1_row4_col2, next_state_share1_row4_col3, next_state_share1_row4_col4 
);
two_dimension_xor inst_next_round_sbox_input_xor_share2 (
add_roundkey_share2_row1_col1, add_roundkey_share2_row1_col2, add_roundkey_share2_row1_col3, add_roundkey_share2_row1_col4, add_roundkey_share2_row2_col1, add_roundkey_share2_row2_col2, add_roundkey_share2_row2_col3, add_roundkey_share2_row2_col4, add_roundkey_share2_row3_col1, add_roundkey_share2_row3_col2, add_roundkey_share2_row3_col3, add_roundkey_share2_row3_col4, add_roundkey_share2_row4_col1, add_roundkey_share2_row4_col2, add_roundkey_share2_row4_col3, add_roundkey_share2_row4_col4 ,
final_sbox_output_share2_row1_col1, final_sbox_output_share2_row1_col2, final_sbox_output_share2_row1_col3, final_sbox_output_share2_row1_col4, final_sbox_output_share2_row2_col1, final_sbox_output_share2_row2_col2, final_sbox_output_share2_row2_col3, final_sbox_output_share2_row2_col4, final_sbox_output_share2_row3_col1, final_sbox_output_share2_row3_col2, final_sbox_output_share2_row3_col3, final_sbox_output_share2_row3_col4, final_sbox_output_share2_row4_col1, final_sbox_output_share2_row4_col2, final_sbox_output_share2_row4_col3, final_sbox_output_share2_row4_col4 ,
next_state_share2_row1_col1, next_state_share2_row1_col2, next_state_share2_row1_col3, next_state_share2_row1_col4, next_state_share2_row2_col1, next_state_share2_row2_col2, next_state_share2_row2_col3, next_state_share2_row2_col4, next_state_share2_row3_col1, next_state_share2_row3_col2, next_state_share2_row3_col3, next_state_share2_row3_col4, next_state_share2_row4_col1, next_state_share2_row4_col2, next_state_share2_row4_col3, next_state_share2_row4_col4 
);

// Control logic
parameter ROUND_STATE_IDLE    = 8'd1 ;
parameter ROUND_STATE_CYCLE1  = 8'd2 ;
parameter ROUND_STATE_CYCLE2  = 8'd3 ;
parameter ROUND_STATE_CYCLE3  = 8'd4 ;
parameter ROUND_STATE_CYCLE4  = 8'd5 ;
parameter ROUND_STATE_CYCLE5  = 8'd6 ;
parameter ROUND_STATE_CYCLE6  = 8'd7 ;
parameter ROUND_STATE_CYCLE7  = 8'd8 ;
parameter ROUND_STATE_CYCLE8  = 8'd9 ;
parameter ROUND_STATE_CYCLE9  = 8'd10;
parameter ROUND_STATE_CYCLE10 = 8'd11;
parameter ROUND_STATE_CYCLE11 = 8'd12;
parameter ROUND_STATE_CYCLE12 = 8'd13;
parameter ROUND_STATE_CYCLE13 = 8'd14;
parameter ROUND_STATE_CYCLE14 = 8'd15;
parameter ROUND_STATE_CYCLE15 = 8'd16;
parameter ROUND_STATE_CYCLE16 = 8'd17;
parameter ROUND_STATE_CYCLE17 = 8'd18;
parameter ROUND_STATE_CYCLE18 = 8'd19;
parameter ROUND_STATE_CYCLE19 = 8'd20;
parameter ROUND_STATE_CYCLE20 = 8'd21;
parameter ROUND_STATE_CYCLE21 = 8'd22;
parameter ROUND_STATE_CYCLE22 = 8'd23;
 
reg [8:1] state_reg, state_next ;
reg in_operation_reg,in_operation_next ;

always@(posedge clk) begin
    if(reset) begin
        state_reg <= ROUND_STATE_IDLE;
        in_operation_reg <= 0;
    end
    else if(start) begin
        state_reg <= ROUND_STATE_CYCLE1;
        in_operation_reg <= 1;
    end
    else begin
        state_reg <= state_next;
        in_operation_reg <= in_operation_next;
    end
end


reg done ;
assign out_done = done;

always@(*) begin
    if(state_reg == ROUND_STATE_IDLE ) begin
        done <= 0;
        state_next <= ROUND_STATE_IDLE;
        in_operation_next <= 0;    
    end
	else if(state_reg == ROUND_STATE_CYCLE21) begin
        done <= 1;
        state_next <= ROUND_STATE_CYCLE21;
        in_operation_next <= 0;    
    end
    else if(in_operation_reg) begin
        done <= 0;
        state_next <= state_reg + 8'd1;
        in_operation_next <= 1;
    end
    else begin
        done <= 0;
        state_next <= state_reg;
		in_operation_next <= in_operation_reg;
    end
end

always@(*) begin
    case (state_reg)
        ROUND_STATE_IDLE: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 1;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 0;    
            select_final_round     <= 0;        
        end
        ROUND_STATE_CYCLE1: begin
            //select_key_state_input <= 1;
            //enable_key_state_input <= 1;
            select_first_round     <= 1;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
        ROUND_STATE_CYCLE2: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end

        ROUND_STATE_CYCLE3: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE4: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end

        ROUND_STATE_CYCLE5: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE6: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end

        ROUND_STATE_CYCLE7: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE8: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end

        ROUND_STATE_CYCLE9: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE10: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end
        ROUND_STATE_CYCLE11: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE12: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end

        ROUND_STATE_CYCLE13: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE14: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end

        ROUND_STATE_CYCLE15: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE16: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end

        ROUND_STATE_CYCLE17: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE18: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 0;        
        end

        ROUND_STATE_CYCLE19: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 1;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 1;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 0;        
        end
		  
        ROUND_STATE_CYCLE20: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 1;            
            select_final_round     <= 1;        
        end

        ROUND_STATE_CYCLE21: begin
            //select_key_state_input <= 0;
            //enable_key_state_input <= 0;
            select_first_round     <= 0;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 0;            
            select_final_round     <= 1;        
        end

        default: begin
            //select_key_state_input <= 1;
            //enable_key_state_input <= 0;
            select_first_round     <= 1;
            enable_sbox_cycle1     <= 0;
            enable_sbox_cycle2     <= 0; 
            select_final_round     <= 0;        
        end
    endcase
end

assign ciphertext_share2 = {next_state_share2_row1_col1, next_state_share2_row2_col1, next_state_share2_row3_col1, next_state_share2_row4_col1, next_state_share2_row1_col2, next_state_share2_row2_col2, next_state_share2_row3_col2, next_state_share2_row4_col2, next_state_share2_row1_col3, next_state_share2_row2_col3, next_state_share2_row3_col3, next_state_share2_row4_col3, next_state_share2_row1_col4, next_state_share2_row2_col4, next_state_share2_row3_col4, next_state_share2_row4_col4 };
assign ciphertext_share1 = {next_state_share1_row1_col1, next_state_share1_row2_col1, next_state_share1_row3_col1, next_state_share1_row4_col1, next_state_share1_row1_col2, next_state_share1_row2_col2, next_state_share1_row3_col2, next_state_share1_row4_col2, next_state_share1_row1_col3, next_state_share1_row2_col3, next_state_share1_row3_col3, next_state_share1_row4_col3, next_state_share1_row1_col4, next_state_share1_row2_col4, next_state_share1_row3_col4, next_state_share1_row4_col4 };

endmodule