`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 02/22/2025
// Design Name: cross_module_multiplication
// Module Name: cross_module_multiplication
// Description: This non-complete module operates on one share from each HO_TSM1 module. 
//              It implements cross multiplication to compute cross-module terms.
// Dependencies: None
// Revision: 0.01 - Initial version
//////////////////////////////////////////////////////////////////////////////////


module cross_module_multiplication (
output_x0_share, output_x1_share, output_x2_share, output_x3_share, output_x0x1_share, output_x0x2_share, output_x0x3_share, output_x1x2_share, output_x1x3_share, output_x2x3_share, output_x0x1x2_share, output_x0x1x3_share, output_x0x2x3_share, output_x1x2x3_share, output_x0x1x2x3_share , 
output_sum_secondmodule_equation_num_0_index_0_share, output_sum_secondmodule_equation_num_0_index_1_share, output_sum_secondmodule_equation_num_0_index_2_share, output_sum_secondmodule_equation_num_0_index_3_share, output_sum_secondmodule_equation_num_0_index_4_share, output_sum_secondmodule_equation_num_0_index_5_share, output_sum_secondmodule_equation_num_0_index_6_share, output_sum_secondmodule_equation_num_0_index_7_share, output_sum_secondmodule_equation_num_0_index_8_share, output_sum_secondmodule_equation_num_0_index_9_share, output_sum_secondmodule_equation_num_0_index_10_share, output_sum_secondmodule_equation_num_0_index_11_share, output_sum_secondmodule_equation_num_0_index_12_share, output_sum_secondmodule_equation_num_0_index_13_share, output_sum_secondmodule_equation_num_0_index_14_share,
output_sum_secondmodule_equation_num_1_index_0_share, output_sum_secondmodule_equation_num_1_index_1_share, output_sum_secondmodule_equation_num_1_index_2_share, output_sum_secondmodule_equation_num_1_index_3_share, output_sum_secondmodule_equation_num_1_index_4_share, output_sum_secondmodule_equation_num_1_index_5_share, output_sum_secondmodule_equation_num_1_index_6_share, output_sum_secondmodule_equation_num_1_index_7_share, output_sum_secondmodule_equation_num_1_index_8_share, output_sum_secondmodule_equation_num_1_index_9_share, output_sum_secondmodule_equation_num_1_index_10_share, output_sum_secondmodule_equation_num_1_index_11_share, output_sum_secondmodule_equation_num_1_index_12_share, output_sum_secondmodule_equation_num_1_index_13_share, output_sum_secondmodule_equation_num_1_index_14_share,
output_sum_secondmodule_equation_num_2_index_0_share, output_sum_secondmodule_equation_num_2_index_1_share, output_sum_secondmodule_equation_num_2_index_2_share, output_sum_secondmodule_equation_num_2_index_3_share, output_sum_secondmodule_equation_num_2_index_4_share, output_sum_secondmodule_equation_num_2_index_5_share, output_sum_secondmodule_equation_num_2_index_6_share, output_sum_secondmodule_equation_num_2_index_7_share, output_sum_secondmodule_equation_num_2_index_8_share, output_sum_secondmodule_equation_num_2_index_9_share, output_sum_secondmodule_equation_num_2_index_10_share, output_sum_secondmodule_equation_num_2_index_11_share, output_sum_secondmodule_equation_num_2_index_12_share, output_sum_secondmodule_equation_num_2_index_13_share, output_sum_secondmodule_equation_num_2_index_14_share,
output_sum_secondmodule_equation_num_3_index_0_share, output_sum_secondmodule_equation_num_3_index_1_share, output_sum_secondmodule_equation_num_3_index_2_share, output_sum_secondmodule_equation_num_3_index_3_share, output_sum_secondmodule_equation_num_3_index_4_share, output_sum_secondmodule_equation_num_3_index_5_share, output_sum_secondmodule_equation_num_3_index_6_share, output_sum_secondmodule_equation_num_3_index_7_share, output_sum_secondmodule_equation_num_3_index_8_share, output_sum_secondmodule_equation_num_3_index_9_share, output_sum_secondmodule_equation_num_3_index_10_share, output_sum_secondmodule_equation_num_3_index_11_share, output_sum_secondmodule_equation_num_3_index_12_share, output_sum_secondmodule_equation_num_3_index_13_share, output_sum_secondmodule_equation_num_3_index_14_share,
output_sum_secondmodule_equation_num_4_index_0_share, output_sum_secondmodule_equation_num_4_index_1_share, output_sum_secondmodule_equation_num_4_index_2_share, output_sum_secondmodule_equation_num_4_index_3_share, output_sum_secondmodule_equation_num_4_index_4_share, output_sum_secondmodule_equation_num_4_index_5_share, output_sum_secondmodule_equation_num_4_index_6_share, output_sum_secondmodule_equation_num_4_index_7_share, output_sum_secondmodule_equation_num_4_index_8_share, output_sum_secondmodule_equation_num_4_index_9_share, output_sum_secondmodule_equation_num_4_index_10_share, output_sum_secondmodule_equation_num_4_index_11_share, output_sum_secondmodule_equation_num_4_index_12_share, output_sum_secondmodule_equation_num_4_index_13_share, output_sum_secondmodule_equation_num_4_index_14_share,
output_sum_secondmodule_equation_num_5_index_0_share, output_sum_secondmodule_equation_num_5_index_1_share, output_sum_secondmodule_equation_num_5_index_2_share, output_sum_secondmodule_equation_num_5_index_3_share, output_sum_secondmodule_equation_num_5_index_4_share, output_sum_secondmodule_equation_num_5_index_5_share, output_sum_secondmodule_equation_num_5_index_6_share, output_sum_secondmodule_equation_num_5_index_7_share, output_sum_secondmodule_equation_num_5_index_8_share, output_sum_secondmodule_equation_num_5_index_9_share, output_sum_secondmodule_equation_num_5_index_10_share, output_sum_secondmodule_equation_num_5_index_11_share, output_sum_secondmodule_equation_num_5_index_12_share, output_sum_secondmodule_equation_num_5_index_13_share, output_sum_secondmodule_equation_num_5_index_14_share,
output_sum_secondmodule_equation_num_6_index_0_share, output_sum_secondmodule_equation_num_6_index_1_share, output_sum_secondmodule_equation_num_6_index_2_share, output_sum_secondmodule_equation_num_6_index_3_share, output_sum_secondmodule_equation_num_6_index_4_share, output_sum_secondmodule_equation_num_6_index_5_share, output_sum_secondmodule_equation_num_6_index_6_share, output_sum_secondmodule_equation_num_6_index_7_share, output_sum_secondmodule_equation_num_6_index_8_share, output_sum_secondmodule_equation_num_6_index_9_share, output_sum_secondmodule_equation_num_6_index_10_share, output_sum_secondmodule_equation_num_6_index_11_share, output_sum_secondmodule_equation_num_6_index_12_share, output_sum_secondmodule_equation_num_6_index_13_share, output_sum_secondmodule_equation_num_6_index_14_share,
output_sum_secondmodule_equation_num_7_index_0_share, output_sum_secondmodule_equation_num_7_index_1_share, output_sum_secondmodule_equation_num_7_index_2_share, output_sum_secondmodule_equation_num_7_index_3_share, output_sum_secondmodule_equation_num_7_index_4_share, output_sum_secondmodule_equation_num_7_index_5_share, output_sum_secondmodule_equation_num_7_index_6_share, output_sum_secondmodule_equation_num_7_index_7_share, output_sum_secondmodule_equation_num_7_index_8_share, output_sum_secondmodule_equation_num_7_index_9_share, output_sum_secondmodule_equation_num_7_index_10_share, output_sum_secondmodule_equation_num_7_index_11_share, output_sum_secondmodule_equation_num_7_index_12_share, output_sum_secondmodule_equation_num_7_index_13_share, output_sum_secondmodule_equation_num_7_index_14_share,
cross_module_equation_num0_domain, cross_module_equation_num1_domain, cross_module_equation_num2_domain, cross_module_equation_num3_domain,cross_module_equation_num4_domain,cross_module_equation_num5_domain,cross_module_equation_num6_domain,cross_module_equation_num7_domain
);

input output_x0_share, output_x1_share, output_x2_share, output_x3_share, output_x0x1_share, output_x0x2_share, output_x0x3_share, output_x1x2_share, output_x1x3_share, output_x2x3_share, output_x0x1x2_share, output_x0x1x3_share, output_x0x2x3_share, output_x1x2x3_share, output_x0x1x2x3_share , 
output_sum_secondmodule_equation_num_0_index_0_share, output_sum_secondmodule_equation_num_0_index_1_share, output_sum_secondmodule_equation_num_0_index_2_share, output_sum_secondmodule_equation_num_0_index_3_share, output_sum_secondmodule_equation_num_0_index_4_share, output_sum_secondmodule_equation_num_0_index_5_share, output_sum_secondmodule_equation_num_0_index_6_share, output_sum_secondmodule_equation_num_0_index_7_share, output_sum_secondmodule_equation_num_0_index_8_share, output_sum_secondmodule_equation_num_0_index_9_share, output_sum_secondmodule_equation_num_0_index_10_share, output_sum_secondmodule_equation_num_0_index_11_share, output_sum_secondmodule_equation_num_0_index_12_share, output_sum_secondmodule_equation_num_0_index_13_share, output_sum_secondmodule_equation_num_0_index_14_share,
output_sum_secondmodule_equation_num_1_index_0_share, output_sum_secondmodule_equation_num_1_index_1_share, output_sum_secondmodule_equation_num_1_index_2_share, output_sum_secondmodule_equation_num_1_index_3_share, output_sum_secondmodule_equation_num_1_index_4_share, output_sum_secondmodule_equation_num_1_index_5_share, output_sum_secondmodule_equation_num_1_index_6_share, output_sum_secondmodule_equation_num_1_index_7_share, output_sum_secondmodule_equation_num_1_index_8_share, output_sum_secondmodule_equation_num_1_index_9_share, output_sum_secondmodule_equation_num_1_index_10_share, output_sum_secondmodule_equation_num_1_index_11_share, output_sum_secondmodule_equation_num_1_index_12_share, output_sum_secondmodule_equation_num_1_index_13_share, output_sum_secondmodule_equation_num_1_index_14_share,
output_sum_secondmodule_equation_num_2_index_0_share, output_sum_secondmodule_equation_num_2_index_1_share, output_sum_secondmodule_equation_num_2_index_2_share, output_sum_secondmodule_equation_num_2_index_3_share, output_sum_secondmodule_equation_num_2_index_4_share, output_sum_secondmodule_equation_num_2_index_5_share, output_sum_secondmodule_equation_num_2_index_6_share, output_sum_secondmodule_equation_num_2_index_7_share, output_sum_secondmodule_equation_num_2_index_8_share, output_sum_secondmodule_equation_num_2_index_9_share, output_sum_secondmodule_equation_num_2_index_10_share, output_sum_secondmodule_equation_num_2_index_11_share, output_sum_secondmodule_equation_num_2_index_12_share, output_sum_secondmodule_equation_num_2_index_13_share, output_sum_secondmodule_equation_num_2_index_14_share,
output_sum_secondmodule_equation_num_3_index_0_share, output_sum_secondmodule_equation_num_3_index_1_share, output_sum_secondmodule_equation_num_3_index_2_share, output_sum_secondmodule_equation_num_3_index_3_share, output_sum_secondmodule_equation_num_3_index_4_share, output_sum_secondmodule_equation_num_3_index_5_share, output_sum_secondmodule_equation_num_3_index_6_share, output_sum_secondmodule_equation_num_3_index_7_share, output_sum_secondmodule_equation_num_3_index_8_share, output_sum_secondmodule_equation_num_3_index_9_share, output_sum_secondmodule_equation_num_3_index_10_share, output_sum_secondmodule_equation_num_3_index_11_share, output_sum_secondmodule_equation_num_3_index_12_share, output_sum_secondmodule_equation_num_3_index_13_share, output_sum_secondmodule_equation_num_3_index_14_share,
output_sum_secondmodule_equation_num_4_index_0_share, output_sum_secondmodule_equation_num_4_index_1_share, output_sum_secondmodule_equation_num_4_index_2_share, output_sum_secondmodule_equation_num_4_index_3_share, output_sum_secondmodule_equation_num_4_index_4_share, output_sum_secondmodule_equation_num_4_index_5_share, output_sum_secondmodule_equation_num_4_index_6_share, output_sum_secondmodule_equation_num_4_index_7_share, output_sum_secondmodule_equation_num_4_index_8_share, output_sum_secondmodule_equation_num_4_index_9_share, output_sum_secondmodule_equation_num_4_index_10_share, output_sum_secondmodule_equation_num_4_index_11_share, output_sum_secondmodule_equation_num_4_index_12_share, output_sum_secondmodule_equation_num_4_index_13_share, output_sum_secondmodule_equation_num_4_index_14_share,
output_sum_secondmodule_equation_num_5_index_0_share, output_sum_secondmodule_equation_num_5_index_1_share, output_sum_secondmodule_equation_num_5_index_2_share, output_sum_secondmodule_equation_num_5_index_3_share, output_sum_secondmodule_equation_num_5_index_4_share, output_sum_secondmodule_equation_num_5_index_5_share, output_sum_secondmodule_equation_num_5_index_6_share, output_sum_secondmodule_equation_num_5_index_7_share, output_sum_secondmodule_equation_num_5_index_8_share, output_sum_secondmodule_equation_num_5_index_9_share, output_sum_secondmodule_equation_num_5_index_10_share, output_sum_secondmodule_equation_num_5_index_11_share, output_sum_secondmodule_equation_num_5_index_12_share, output_sum_secondmodule_equation_num_5_index_13_share, output_sum_secondmodule_equation_num_5_index_14_share,
output_sum_secondmodule_equation_num_6_index_0_share, output_sum_secondmodule_equation_num_6_index_1_share, output_sum_secondmodule_equation_num_6_index_2_share, output_sum_secondmodule_equation_num_6_index_3_share, output_sum_secondmodule_equation_num_6_index_4_share, output_sum_secondmodule_equation_num_6_index_5_share, output_sum_secondmodule_equation_num_6_index_6_share, output_sum_secondmodule_equation_num_6_index_7_share, output_sum_secondmodule_equation_num_6_index_8_share, output_sum_secondmodule_equation_num_6_index_9_share, output_sum_secondmodule_equation_num_6_index_10_share, output_sum_secondmodule_equation_num_6_index_11_share, output_sum_secondmodule_equation_num_6_index_12_share, output_sum_secondmodule_equation_num_6_index_13_share, output_sum_secondmodule_equation_num_6_index_14_share,
output_sum_secondmodule_equation_num_7_index_0_share, output_sum_secondmodule_equation_num_7_index_1_share, output_sum_secondmodule_equation_num_7_index_2_share, output_sum_secondmodule_equation_num_7_index_3_share, output_sum_secondmodule_equation_num_7_index_4_share, output_sum_secondmodule_equation_num_7_index_5_share, output_sum_secondmodule_equation_num_7_index_6_share, output_sum_secondmodule_equation_num_7_index_7_share, output_sum_secondmodule_equation_num_7_index_8_share, output_sum_secondmodule_equation_num_7_index_9_share, output_sum_secondmodule_equation_num_7_index_10_share, output_sum_secondmodule_equation_num_7_index_11_share, output_sum_secondmodule_equation_num_7_index_12_share, output_sum_secondmodule_equation_num_7_index_13_share, output_sum_secondmodule_equation_num_7_index_14_share;

output cross_module_equation_num0_domain, cross_module_equation_num1_domain, cross_module_equation_num2_domain, cross_module_equation_num3_domain,cross_module_equation_num4_domain,cross_module_equation_num5_domain,cross_module_equation_num6_domain,cross_module_equation_num7_domain ;



assign cross_module_equation_num0_domain = output_x0_share &output_sum_secondmodule_equation_num_0_index_0_share ^  output_x1_share &output_sum_secondmodule_equation_num_0_index_1_share ^  output_x2_share &output_sum_secondmodule_equation_num_0_index_2_share ^  output_x3_share &output_sum_secondmodule_equation_num_0_index_3_share ^  output_x0x1_share &output_sum_secondmodule_equation_num_0_index_4_share ^  output_x0x2_share &output_sum_secondmodule_equation_num_0_index_5_share ^  output_x0x3_share &output_sum_secondmodule_equation_num_0_index_6_share ^  output_x1x2_share &output_sum_secondmodule_equation_num_0_index_7_share ^  output_x1x3_share &output_sum_secondmodule_equation_num_0_index_8_share ^  output_x2x3_share &output_sum_secondmodule_equation_num_0_index_9_share ^  output_x0x1x2_share &output_sum_secondmodule_equation_num_0_index_10_share ^  output_x0x1x3_share &output_sum_secondmodule_equation_num_0_index_11_share ^  output_x0x2x3_share &output_sum_secondmodule_equation_num_0_index_12_share ^  output_x1x2x3_share &output_sum_secondmodule_equation_num_0_index_13_share ^  output_x0x1x2x3_share &output_sum_secondmodule_equation_num_0_index_14_share  ;
assign cross_module_equation_num1_domain = output_x0_share &output_sum_secondmodule_equation_num_1_index_0_share ^  output_x1_share &output_sum_secondmodule_equation_num_1_index_1_share ^  output_x2_share &output_sum_secondmodule_equation_num_1_index_2_share ^  output_x3_share &output_sum_secondmodule_equation_num_1_index_3_share ^  output_x0x1_share &output_sum_secondmodule_equation_num_1_index_4_share ^  output_x0x2_share &output_sum_secondmodule_equation_num_1_index_5_share ^  output_x0x3_share &output_sum_secondmodule_equation_num_1_index_6_share ^  output_x1x2_share &output_sum_secondmodule_equation_num_1_index_7_share ^  output_x1x3_share &output_sum_secondmodule_equation_num_1_index_8_share ^  output_x2x3_share &output_sum_secondmodule_equation_num_1_index_9_share ^  output_x0x1x2_share &output_sum_secondmodule_equation_num_1_index_10_share ^  output_x0x1x3_share &output_sum_secondmodule_equation_num_1_index_11_share ^  output_x0x2x3_share &output_sum_secondmodule_equation_num_1_index_12_share ^  output_x1x2x3_share &output_sum_secondmodule_equation_num_1_index_13_share ^  output_x0x1x2x3_share &output_sum_secondmodule_equation_num_1_index_14_share  ;
assign cross_module_equation_num2_domain = output_x0_share &output_sum_secondmodule_equation_num_2_index_0_share ^  output_x1_share &output_sum_secondmodule_equation_num_2_index_1_share ^  output_x2_share &output_sum_secondmodule_equation_num_2_index_2_share ^  output_x3_share &output_sum_secondmodule_equation_num_2_index_3_share ^  output_x0x1_share &output_sum_secondmodule_equation_num_2_index_4_share ^  output_x0x2_share &output_sum_secondmodule_equation_num_2_index_5_share ^  output_x0x3_share &output_sum_secondmodule_equation_num_2_index_6_share ^  output_x1x2_share &output_sum_secondmodule_equation_num_2_index_7_share ^  output_x1x3_share &output_sum_secondmodule_equation_num_2_index_8_share ^  output_x2x3_share &output_sum_secondmodule_equation_num_2_index_9_share ^  output_x0x1x2_share &output_sum_secondmodule_equation_num_2_index_10_share ^  output_x0x1x3_share &output_sum_secondmodule_equation_num_2_index_11_share ^  output_x0x2x3_share &output_sum_secondmodule_equation_num_2_index_12_share ^  output_x1x2x3_share &output_sum_secondmodule_equation_num_2_index_13_share ^  output_x0x1x2x3_share &output_sum_secondmodule_equation_num_2_index_14_share  ;
assign cross_module_equation_num3_domain = output_x0_share &output_sum_secondmodule_equation_num_3_index_0_share ^  output_x1_share &output_sum_secondmodule_equation_num_3_index_1_share ^  output_x2_share &output_sum_secondmodule_equation_num_3_index_2_share ^  output_x3_share &output_sum_secondmodule_equation_num_3_index_3_share ^  output_x0x1_share &output_sum_secondmodule_equation_num_3_index_4_share ^  output_x0x2_share &output_sum_secondmodule_equation_num_3_index_5_share ^  output_x0x3_share &output_sum_secondmodule_equation_num_3_index_6_share ^  output_x1x2_share &output_sum_secondmodule_equation_num_3_index_7_share ^  output_x1x3_share &output_sum_secondmodule_equation_num_3_index_8_share ^  output_x2x3_share &output_sum_secondmodule_equation_num_3_index_9_share ^  output_x0x1x2_share &output_sum_secondmodule_equation_num_3_index_10_share ^  output_x0x1x3_share &output_sum_secondmodule_equation_num_3_index_11_share ^  output_x0x2x3_share &output_sum_secondmodule_equation_num_3_index_12_share ^  output_x1x2x3_share &output_sum_secondmodule_equation_num_3_index_13_share ^  output_x0x1x2x3_share &output_sum_secondmodule_equation_num_3_index_14_share  ;
assign cross_module_equation_num4_domain = output_x0_share &output_sum_secondmodule_equation_num_4_index_0_share ^  output_x1_share &output_sum_secondmodule_equation_num_4_index_1_share ^  output_x2_share &output_sum_secondmodule_equation_num_4_index_2_share ^  output_x3_share &output_sum_secondmodule_equation_num_4_index_3_share ^  output_x0x1_share &output_sum_secondmodule_equation_num_4_index_4_share ^  output_x0x2_share &output_sum_secondmodule_equation_num_4_index_5_share ^  output_x0x3_share &output_sum_secondmodule_equation_num_4_index_6_share ^  output_x1x2_share &output_sum_secondmodule_equation_num_4_index_7_share ^  output_x1x3_share &output_sum_secondmodule_equation_num_4_index_8_share ^  output_x2x3_share &output_sum_secondmodule_equation_num_4_index_9_share ^  output_x0x1x2_share &output_sum_secondmodule_equation_num_4_index_10_share ^  output_x0x1x3_share &output_sum_secondmodule_equation_num_4_index_11_share ^  output_x0x2x3_share &output_sum_secondmodule_equation_num_4_index_12_share ^  output_x1x2x3_share &output_sum_secondmodule_equation_num_4_index_13_share ^  output_x0x1x2x3_share &output_sum_secondmodule_equation_num_4_index_14_share  ;
assign cross_module_equation_num5_domain = output_x0_share &output_sum_secondmodule_equation_num_5_index_0_share ^  output_x1_share &output_sum_secondmodule_equation_num_5_index_1_share ^  output_x2_share &output_sum_secondmodule_equation_num_5_index_2_share ^  output_x3_share &output_sum_secondmodule_equation_num_5_index_3_share ^  output_x0x1_share &output_sum_secondmodule_equation_num_5_index_4_share ^  output_x0x2_share &output_sum_secondmodule_equation_num_5_index_5_share ^  output_x0x3_share &output_sum_secondmodule_equation_num_5_index_6_share ^  output_x1x2_share &output_sum_secondmodule_equation_num_5_index_7_share ^  output_x1x3_share &output_sum_secondmodule_equation_num_5_index_8_share ^  output_x2x3_share &output_sum_secondmodule_equation_num_5_index_9_share ^  output_x0x1x2_share &output_sum_secondmodule_equation_num_5_index_10_share ^  output_x0x1x3_share &output_sum_secondmodule_equation_num_5_index_11_share ^  output_x0x2x3_share &output_sum_secondmodule_equation_num_5_index_12_share ^  output_x1x2x3_share &output_sum_secondmodule_equation_num_5_index_13_share ^  output_x0x1x2x3_share &output_sum_secondmodule_equation_num_5_index_14_share  ;
assign cross_module_equation_num6_domain = output_x0_share &output_sum_secondmodule_equation_num_6_index_0_share ^  output_x1_share &output_sum_secondmodule_equation_num_6_index_1_share ^  output_x2_share &output_sum_secondmodule_equation_num_6_index_2_share ^  output_x3_share &output_sum_secondmodule_equation_num_6_index_3_share ^  output_x0x1_share &output_sum_secondmodule_equation_num_6_index_4_share ^  output_x0x2_share &output_sum_secondmodule_equation_num_6_index_5_share ^  output_x0x3_share &output_sum_secondmodule_equation_num_6_index_6_share ^  output_x1x2_share &output_sum_secondmodule_equation_num_6_index_7_share ^  output_x1x3_share &output_sum_secondmodule_equation_num_6_index_8_share ^  output_x2x3_share &output_sum_secondmodule_equation_num_6_index_9_share ^  output_x0x1x2_share &output_sum_secondmodule_equation_num_6_index_10_share ^  output_x0x1x3_share &output_sum_secondmodule_equation_num_6_index_11_share ^  output_x0x2x3_share &output_sum_secondmodule_equation_num_6_index_12_share ^  output_x1x2x3_share &output_sum_secondmodule_equation_num_6_index_13_share ^  output_x0x1x2x3_share &output_sum_secondmodule_equation_num_6_index_14_share  ;
assign cross_module_equation_num7_domain = output_x0_share &output_sum_secondmodule_equation_num_7_index_0_share ^  output_x1_share &output_sum_secondmodule_equation_num_7_index_1_share ^  output_x2_share &output_sum_secondmodule_equation_num_7_index_2_share ^  output_x3_share &output_sum_secondmodule_equation_num_7_index_3_share ^  output_x0x1_share &output_sum_secondmodule_equation_num_7_index_4_share ^  output_x0x2_share &output_sum_secondmodule_equation_num_7_index_5_share ^  output_x0x3_share &output_sum_secondmodule_equation_num_7_index_6_share ^  output_x1x2_share &output_sum_secondmodule_equation_num_7_index_7_share ^  output_x1x3_share &output_sum_secondmodule_equation_num_7_index_8_share ^  output_x2x3_share &output_sum_secondmodule_equation_num_7_index_9_share ^  output_x0x1x2_share &output_sum_secondmodule_equation_num_7_index_10_share ^  output_x0x1x3_share &output_sum_secondmodule_equation_num_7_index_11_share ^  output_x0x2x3_share &output_sum_secondmodule_equation_num_7_index_12_share ^  output_x1x2x3_share &output_sum_secondmodule_equation_num_7_index_13_share ^  output_x0x1x2x3_share &output_sum_secondmodule_equation_num_7_index_14_share  ;


endmodule