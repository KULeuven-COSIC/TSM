`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 22:00:00 02/22/2025
// Design Name: All Cross Products of One Share
// Module Name: allcrossproducts_oneshare_eightinputs
// Project Name: AES Masked S-Box
// Description: Computes all cross-products of 8 inputs for exactly one share.
// Dependencies: None
//
// Revision:
// Revision 0.01 - File Created
//
//////////////////////////////////////////////////////////////////////////////////

module allcrossproducts_oneshare_eightinputs(
x0_share_in, x1_share_in, x2_share_in, x3_share_in, x4_share_in, x5_share_in, x6_share_in, x7_share_in ,
x0_share_out             , x1_share_out             , x2_share_out             , x3_share_out             , x4_share_out             , x5_share_out             , x6_share_out             , x7_share_out             , x0x1_share_out           , x0x4_share_out           , x0x5_share_out           , x0x6_share_out           , x1x2_share_out           , x1x3_share_out           , x1x4_share_out           , x1x6_share_out           , x2x3_share_out           , x2x4_share_out           , x2x6_share_out           , x2x7_share_out           , x4x6_share_out           , x5x6_share_out           , x5x7_share_out           , x6x7_share_out           , x0x2_share_out           , x0x3_share_out           , x0x7_share_out           , x1x7_share_out           , x3x7_share_out           , x4x5_share_out           , x3x4_share_out           , x4x7_share_out           , x3x6_share_out           , x1x5_share_out           , x2x5_share_out           , x3x5_share_out           , x0x1x4_share_out         , x0x1x6_share_out         , x0x1x7_share_out         , x0x2x4_share_out         , x0x2x5_share_out         , x0x2x6_share_out         , x0x2x7_share_out         , x0x3x4_share_out         , x0x3x5_share_out         , x0x3x6_share_out         , x0x4x6_share_out         , x0x4x7_share_out         , x1x2x3_share_out         , x1x2x4_share_out         , x1x2x6_share_out         , x1x3x4_share_out         , x1x3x7_share_out         , x1x4x6_share_out         , x1x5x6_share_out         , x2x3x5_share_out         , x2x3x7_share_out         , x2x4x7_share_out         , x2x5x6_share_out         , x2x5x7_share_out         , x2x6x7_share_out         , x3x4x7_share_out         , x3x5x7_share_out         , x3x6x7_share_out         , x4x5x6_share_out         , x5x6x7_share_out         , x0x1x3_share_out         , x0x2x3_share_out         , x0x4x5_share_out         , x0x5x7_share_out         , x0x6x7_share_out         , x1x3x5_share_out         , x1x3x6_share_out         , x1x4x7_share_out         , x2x3x4_share_out         , x2x3x6_share_out         , x3x4x6_share_out         , x3x5x6_share_out         , x0x1x5_share_out         , x0x3x7_share_out         , x1x2x5_share_out         , x1x2x7_share_out         , x1x4x5_share_out         , x1x5x7_share_out         , x2x4x5_share_out         , x3x4x5_share_out         , x4x6x7_share_out         , x1x6x7_share_out         , x4x5x7_share_out         , x0x1x2_share_out         , x0x5x6_share_out         , x2x4x6_share_out         , x0x1x2x3_share_out       , x0x1x2x5_share_out       , x0x1x2x6_share_out       , x0x1x2x7_share_out       , x0x1x4x5_share_out       , x0x1x4x7_share_out       , x0x2x3x5_share_out       , x0x2x3x7_share_out       , x0x2x4x5_share_out       , x0x2x4x7_share_out       , x0x2x5x6_share_out       , x0x2x5x7_share_out       , x0x3x4x6_share_out       , x0x3x5x6_share_out       , x0x4x5x6_share_out       , x0x4x5x7_share_out       , x0x4x6x7_share_out       , x1x2x3x5_share_out       , x1x2x3x6_share_out       , x1x2x3x7_share_out       , x1x2x4x6_share_out       , x1x2x4x7_share_out       , x1x2x6x7_share_out       , x1x3x4x6_share_out       , x1x3x6x7_share_out       , x1x4x5x6_share_out       , x1x4x5x7_share_out       , x1x5x6x7_share_out       , x2x3x5x7_share_out       , x2x3x6x7_share_out       , x2x4x5x6_share_out       , x2x4x5x7_share_out       , x3x5x6x7_share_out       , x0x1x3x4_share_out       , x0x1x3x6_share_out       , x0x1x5x6_share_out       , x0x2x3x6_share_out       , x0x3x4x5_share_out       , x1x2x5x6_share_out       , x1x2x5x7_share_out       , x1x3x4x5_share_out       , x1x3x4x7_share_out       , x1x3x5x6_share_out       , x1x3x5x7_share_out       , x1x4x6x7_share_out       , x2x3x4x5_share_out       , x2x3x4x7_share_out       , x2x4x6x7_share_out       , x3x4x5x6_share_out       , x3x4x5x7_share_out       , x3x4x6x7_share_out       , x0x1x3x5_share_out       , x0x1x4x6_share_out       , x0x2x3x4_share_out       , x0x2x4x6_share_out       , x0x3x4x7_share_out       , x0x3x5x7_share_out       , x1x2x3x4_share_out       , x2x3x4x6_share_out       , x2x3x5x6_share_out       , x2x5x6x7_share_out       , x4x5x6x7_share_out       , x0x1x2x4_share_out       , x0x1x6x7_share_out       , x0x2x6x7_share_out       , x0x3x6x7_share_out       , x0x5x6x7_share_out       , x1x2x4x5_share_out       , x0x1x3x7_share_out       , x0x1x5x7_share_out       , x0x1x2x3x4_share_out     , x0x1x2x3x6_share_out     , x0x1x2x3x7_share_out     , x0x1x2x4x5_share_out     , x0x1x2x4x7_share_out     , x0x1x2x5x7_share_out     , x0x1x2x6x7_share_out     , x0x1x3x4x6_share_out     , x0x1x3x5x6_share_out     , x0x1x3x5x7_share_out     , x0x1x3x6x7_share_out     , x0x1x4x5x6_share_out     , x0x1x5x6x7_share_out     , x0x2x3x4x5_share_out     , x0x2x3x4x6_share_out     , x0x2x4x5x7_share_out     , x0x2x4x6x7_share_out     , x0x3x4x5x6_share_out     , x0x3x4x5x7_share_out     , x0x3x4x6x7_share_out     , x0x3x5x6x7_share_out     , x1x2x3x5x6_share_out     , x1x2x3x5x7_share_out     , x1x2x4x5x6_share_out     , x1x2x4x6x7_share_out     , x1x2x5x6x7_share_out     , x1x3x4x5x7_share_out     , x2x3x4x5x6_share_out     , x2x3x4x5x7_share_out     , x2x4x5x6x7_share_out     , x0x1x2x4x6_share_out     , x0x1x3x4x7_share_out     , x0x2x3x4x7_share_out     , x0x2x3x5x7_share_out     , x0x2x3x6x7_share_out     , x0x2x4x5x6_share_out     , x0x2x5x6x7_share_out     , x0x4x5x6x7_share_out     , x1x2x3x4x6_share_out     , x1x3x4x5x6_share_out     , x2x3x4x6x7_share_out     , x0x1x2x3x5_share_out     , x0x1x4x6x7_share_out     , x1x2x3x4x5_share_out     , x1x2x3x6x7_share_out     , x1x2x4x5x7_share_out     , x1x3x4x6x7_share_out     , x1x3x5x6x7_share_out     , x1x4x5x6x7_share_out     , x2x3x5x6x7_share_out     , x3x4x5x6x7_share_out     , x0x1x2x5x6_share_out     , x0x1x3x4x5_share_out     , x0x1x4x5x7_share_out     , x0x2x3x5x6_share_out     , x1x2x3x4x7_share_out     , x0x1x2x3x4x6_share_out   , x0x1x2x3x4x7_share_out   , x0x1x2x3x5x7_share_out   , x0x1x2x3x6x7_share_out   , x0x1x2x4x5x7_share_out   , x0x1x2x5x6x7_share_out   , x0x1x3x4x6x7_share_out   , x0x1x4x5x6x7_share_out   , x0x2x3x4x5x6_share_out   , x0x2x3x4x5x7_share_out   , x0x2x3x5x6x7_share_out   , x1x2x3x4x6x7_share_out   , x1x2x4x5x6x7_share_out   , x1x3x4x5x6x7_share_out   , x2x3x4x5x6x7_share_out   , x0x1x2x3x5x6_share_out   , x0x1x2x4x6x7_share_out   , x0x1x3x4x5x6_share_out   , x0x2x3x4x6x7_share_out   , x1x2x3x4x5x6_share_out   , x1x2x3x5x6x7_share_out   , x0x1x2x3x4x5_share_out   , x0x1x2x4x5x6_share_out   , x0x1x3x4x5x7_share_out   , x0x1x3x5x6x7_share_out   , x0x2x4x5x6x7_share_out   , x1x2x3x4x5x7_share_out   , x0x3x4x5x6x7_share_out   , x0x1x2x3x4x6x7_share_out , x0x1x2x4x5x6x7_share_out , x0x2x3x4x5x6x7_share_out , x0x1x2x3x5x6x7_share_out , x0x1x3x4x5x6x7_share_out , x1x2x3x4x5x6x7_share_out , x0x1x2x3x4x5x6_share_out , x0x1x2x3x4x5x7_share_out
);

input  x0_share_in, x1_share_in, x2_share_in, x3_share_in, x4_share_in, x5_share_in, x6_share_in, x7_share_in ;
output x0_share_out             , x1_share_out             , x2_share_out             , x3_share_out             , x4_share_out             , x5_share_out             , x6_share_out             , x7_share_out             , x0x1_share_out           , x0x4_share_out           , x0x5_share_out           , x0x6_share_out           , x1x2_share_out           , x1x3_share_out           , x1x4_share_out           , x1x6_share_out           , x2x3_share_out           , x2x4_share_out           , x2x6_share_out           , x2x7_share_out           , x4x6_share_out           , x5x6_share_out           , x5x7_share_out           , x6x7_share_out           , x0x2_share_out           , x0x3_share_out           , x0x7_share_out           , x1x7_share_out           , x3x7_share_out           , x4x5_share_out           , x3x4_share_out           , x4x7_share_out           , x3x6_share_out           , x1x5_share_out           , x2x5_share_out           , x3x5_share_out           , x0x1x4_share_out         , x0x1x6_share_out         , x0x1x7_share_out         , x0x2x4_share_out         , x0x2x5_share_out         , x0x2x6_share_out         , x0x2x7_share_out         , x0x3x4_share_out         , x0x3x5_share_out         , x0x3x6_share_out         , x0x4x6_share_out         , x0x4x7_share_out         , x1x2x3_share_out         , x1x2x4_share_out         , x1x2x6_share_out         , x1x3x4_share_out         , x1x3x7_share_out         , x1x4x6_share_out         , x1x5x6_share_out         , x2x3x5_share_out         , x2x3x7_share_out         , x2x4x7_share_out         , x2x5x6_share_out         , x2x5x7_share_out         , x2x6x7_share_out         , x3x4x7_share_out         , x3x5x7_share_out         , x3x6x7_share_out         , x4x5x6_share_out         , x5x6x7_share_out         , x0x1x3_share_out         , x0x2x3_share_out         , x0x4x5_share_out         , x0x5x7_share_out         , x0x6x7_share_out         , x1x3x5_share_out         , x1x3x6_share_out         , x1x4x7_share_out         , x2x3x4_share_out         , x2x3x6_share_out         , x3x4x6_share_out         , x3x5x6_share_out         , x0x1x5_share_out         , x0x3x7_share_out         , x1x2x5_share_out         , x1x2x7_share_out         , x1x4x5_share_out         , x1x5x7_share_out         , x2x4x5_share_out         , x3x4x5_share_out         , x4x6x7_share_out         , x1x6x7_share_out         , x4x5x7_share_out         , x0x1x2_share_out         , x0x5x6_share_out         , x2x4x6_share_out         , x0x1x2x3_share_out       , x0x1x2x5_share_out       , x0x1x2x6_share_out       , x0x1x2x7_share_out       , x0x1x4x5_share_out       , x0x1x4x7_share_out       , x0x2x3x5_share_out       , x0x2x3x7_share_out       , x0x2x4x5_share_out       , x0x2x4x7_share_out       , x0x2x5x6_share_out       , x0x2x5x7_share_out       , x0x3x4x6_share_out       , x0x3x5x6_share_out       , x0x4x5x6_share_out       , x0x4x5x7_share_out       , x0x4x6x7_share_out       , x1x2x3x5_share_out       , x1x2x3x6_share_out       , x1x2x3x7_share_out       , x1x2x4x6_share_out       , x1x2x4x7_share_out       , x1x2x6x7_share_out       , x1x3x4x6_share_out       , x1x3x6x7_share_out       , x1x4x5x6_share_out       , x1x4x5x7_share_out       , x1x5x6x7_share_out       , x2x3x5x7_share_out       , x2x3x6x7_share_out       , x2x4x5x6_share_out       , x2x4x5x7_share_out       , x3x5x6x7_share_out       , x0x1x3x4_share_out       , x0x1x3x6_share_out       , x0x1x5x6_share_out       , x0x2x3x6_share_out       , x0x3x4x5_share_out       , x1x2x5x6_share_out       , x1x2x5x7_share_out       , x1x3x4x5_share_out       , x1x3x4x7_share_out       , x1x3x5x6_share_out       , x1x3x5x7_share_out       , x1x4x6x7_share_out       , x2x3x4x5_share_out       , x2x3x4x7_share_out       , x2x4x6x7_share_out       , x3x4x5x6_share_out       , x3x4x5x7_share_out       , x3x4x6x7_share_out       , x0x1x3x5_share_out       , x0x1x4x6_share_out       , x0x2x3x4_share_out       , x0x2x4x6_share_out       , x0x3x4x7_share_out       , x0x3x5x7_share_out       , x1x2x3x4_share_out       , x2x3x4x6_share_out       , x2x3x5x6_share_out       , x2x5x6x7_share_out       , x4x5x6x7_share_out       , x0x1x2x4_share_out       , x0x1x6x7_share_out       , x0x2x6x7_share_out       , x0x3x6x7_share_out       , x0x5x6x7_share_out       , x1x2x4x5_share_out       , x0x1x3x7_share_out       , x0x1x5x7_share_out       , x0x1x2x3x4_share_out     , x0x1x2x3x6_share_out     , x0x1x2x3x7_share_out     , x0x1x2x4x5_share_out     , x0x1x2x4x7_share_out     , x0x1x2x5x7_share_out     , x0x1x2x6x7_share_out     , x0x1x3x4x6_share_out     , x0x1x3x5x6_share_out     , x0x1x3x5x7_share_out     , x0x1x3x6x7_share_out     , x0x1x4x5x6_share_out     , x0x1x5x6x7_share_out     , x0x2x3x4x5_share_out     , x0x2x3x4x6_share_out     , x0x2x4x5x7_share_out     , x0x2x4x6x7_share_out     , x0x3x4x5x6_share_out     , x0x3x4x5x7_share_out     , x0x3x4x6x7_share_out     , x0x3x5x6x7_share_out     , x1x2x3x5x6_share_out     , x1x2x3x5x7_share_out     , x1x2x4x5x6_share_out     , x1x2x4x6x7_share_out     , x1x2x5x6x7_share_out     , x1x3x4x5x7_share_out     , x2x3x4x5x6_share_out     , x2x3x4x5x7_share_out     , x2x4x5x6x7_share_out     , x0x1x2x4x6_share_out     , x0x1x3x4x7_share_out     , x0x2x3x4x7_share_out     , x0x2x3x5x7_share_out     , x0x2x3x6x7_share_out     , x0x2x4x5x6_share_out     , x0x2x5x6x7_share_out     , x0x4x5x6x7_share_out     , x1x2x3x4x6_share_out     , x1x3x4x5x6_share_out     , x2x3x4x6x7_share_out     , x0x1x2x3x5_share_out     , x0x1x4x6x7_share_out     , x1x2x3x4x5_share_out     , x1x2x3x6x7_share_out     , x1x2x4x5x7_share_out     , x1x3x4x6x7_share_out     , x1x3x5x6x7_share_out     , x1x4x5x6x7_share_out     , x2x3x5x6x7_share_out     , x3x4x5x6x7_share_out     , x0x1x2x5x6_share_out     , x0x1x3x4x5_share_out     , x0x1x4x5x7_share_out     , x0x2x3x5x6_share_out     , x1x2x3x4x7_share_out     , x0x1x2x3x4x6_share_out   , x0x1x2x3x4x7_share_out   , x0x1x2x3x5x7_share_out   , x0x1x2x3x6x7_share_out   , x0x1x2x4x5x7_share_out   , x0x1x2x5x6x7_share_out   , x0x1x3x4x6x7_share_out   , x0x1x4x5x6x7_share_out   , x0x2x3x4x5x6_share_out   , x0x2x3x4x5x7_share_out   , x0x2x3x5x6x7_share_out   , x1x2x3x4x6x7_share_out   , x1x2x4x5x6x7_share_out   , x1x3x4x5x6x7_share_out   , x2x3x4x5x6x7_share_out   , x0x1x2x3x5x6_share_out   , x0x1x2x4x6x7_share_out   , x0x1x3x4x5x6_share_out   , x0x2x3x4x6x7_share_out   , x1x2x3x4x5x6_share_out   , x1x2x3x5x6x7_share_out   , x0x1x2x3x4x5_share_out   , x0x1x2x4x5x6_share_out   , x0x1x3x4x5x7_share_out   , x0x1x3x5x6x7_share_out   , x0x2x4x5x6x7_share_out   , x1x2x3x4x5x7_share_out   , x0x3x4x5x6x7_share_out   , x0x1x2x3x4x6x7_share_out , x0x1x2x4x5x6x7_share_out , x0x2x3x4x5x6x7_share_out , x0x1x2x3x5x6x7_share_out , x0x1x3x4x5x6x7_share_out , x1x2x3x4x5x6x7_share_out , x0x1x2x3x4x5x6_share_out , x0x1x2x3x4x5x7_share_out ;

assign x0_share_out             =  x0_share_in ;
assign x1_share_out             =  x1_share_in ;
assign x2_share_out             =  x2_share_in ;
assign x3_share_out             =  x3_share_in ;
assign x4_share_out             =  x4_share_in ;
assign x5_share_out             =  x5_share_in ;
assign x6_share_out             =  x6_share_in ;
assign x7_share_out             =  x7_share_in ;
assign x0x1_share_out           =  x0_share_in & x1_share_in   ;
assign x0x4_share_out           =  x0_share_in & x4_share_in   ;
assign x0x5_share_out           =  x0_share_in & x5_share_in   ;
assign x0x6_share_out           =  x0_share_in & x6_share_in   ;
assign x1x2_share_out           =  x1_share_in & x2_share_in   ;
assign x1x3_share_out           =  x1_share_in & x3_share_in   ;
assign x1x4_share_out           =  x1_share_in & x4_share_in   ;
assign x1x6_share_out           =  x1_share_in & x6_share_in   ;
assign x2x3_share_out           =  x2_share_in & x3_share_in   ;
assign x2x4_share_out           =  x2_share_in & x4_share_in   ;
assign x2x6_share_out           =  x2_share_in & x6_share_in   ;
assign x2x7_share_out           =  x2_share_in & x7_share_in   ;
assign x4x6_share_out           =  x4_share_in & x6_share_in   ;
assign x5x6_share_out           =  x5_share_in & x6_share_in   ;
assign x5x7_share_out           =  x5_share_in & x7_share_in   ;
assign x6x7_share_out           =  x6_share_in & x7_share_in   ;
assign x0x2_share_out           =  x0_share_in & x2_share_in   ;
assign x0x3_share_out           =  x0_share_in & x3_share_in   ;
assign x0x7_share_out           =  x0_share_in & x7_share_in   ;
assign x1x7_share_out           =  x1_share_in & x7_share_in   ;
assign x3x7_share_out           =  x3_share_in & x7_share_in   ;
assign x4x5_share_out           =  x4_share_in & x5_share_in   ;
assign x3x4_share_out           =  x3_share_in & x4_share_in   ;
assign x4x7_share_out           =  x4_share_in & x7_share_in   ;
assign x3x6_share_out           =  x3_share_in & x6_share_in   ;
assign x1x5_share_out           =  x1_share_in & x5_share_in   ;
assign x2x5_share_out           =  x2_share_in & x5_share_in   ;
assign x3x5_share_out           =  x3_share_in & x5_share_in   ;
assign x0x1x4_share_out         =  x0_share_in & x1_share_in & x4_share_in   ;
assign x0x1x6_share_out         =  x0_share_in & x1_share_in & x6_share_in   ;
assign x0x1x7_share_out         =  x0_share_in & x1_share_in & x7_share_in   ;
assign x0x2x4_share_out         =  x0_share_in & x2_share_in & x4_share_in   ;
assign x0x2x5_share_out         =  x0_share_in & x2_share_in & x5_share_in   ;
assign x0x2x6_share_out         =  x0_share_in & x2_share_in & x6_share_in   ;
assign x0x2x7_share_out         =  x0_share_in & x2_share_in & x7_share_in   ;
assign x0x3x4_share_out         =  x0_share_in & x3_share_in & x4_share_in   ;
assign x0x3x5_share_out         =  x0_share_in & x3_share_in & x5_share_in   ;
assign x0x3x6_share_out         =  x0_share_in & x3_share_in & x6_share_in   ;
assign x0x4x6_share_out         =  x0_share_in & x4_share_in & x6_share_in   ;
assign x0x4x7_share_out         =  x0_share_in & x4_share_in & x7_share_in   ;
assign x1x2x3_share_out         =  x1_share_in & x2_share_in & x3_share_in   ;
assign x1x2x4_share_out         =  x1_share_in & x2_share_in & x4_share_in   ;
assign x1x2x6_share_out         =  x1_share_in & x2_share_in & x6_share_in   ;
assign x1x3x4_share_out         =  x1_share_in & x3_share_in & x4_share_in   ;
assign x1x3x7_share_out         =  x1_share_in & x3_share_in & x7_share_in   ;
assign x1x4x6_share_out         =  x1_share_in & x4_share_in & x6_share_in   ;
assign x1x5x6_share_out         =  x1_share_in & x5_share_in & x6_share_in   ;
assign x2x3x5_share_out         =  x2_share_in & x3_share_in & x5_share_in   ;
assign x2x3x7_share_out         =  x2_share_in & x3_share_in & x7_share_in   ;
assign x2x4x7_share_out         =  x2_share_in & x4_share_in & x7_share_in   ;
assign x2x5x6_share_out         =  x2_share_in & x5_share_in & x6_share_in   ;
assign x2x5x7_share_out         =  x2_share_in & x5_share_in & x7_share_in   ;
assign x2x6x7_share_out         =  x2_share_in & x6_share_in & x7_share_in   ;
assign x3x4x7_share_out         =  x3_share_in & x4_share_in & x7_share_in   ;
assign x3x5x7_share_out         =  x3_share_in & x5_share_in & x7_share_in   ;
assign x3x6x7_share_out         =  x3_share_in & x6_share_in & x7_share_in   ;
assign x4x5x6_share_out         =  x4_share_in & x5_share_in & x6_share_in   ;
assign x5x6x7_share_out         =  x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3_share_out         =  x0_share_in & x1_share_in & x3_share_in   ;
assign x0x2x3_share_out         =  x0_share_in & x2_share_in & x3_share_in   ;
assign x0x4x5_share_out         =  x0_share_in & x4_share_in & x5_share_in   ;
assign x0x5x7_share_out         =  x0_share_in & x5_share_in & x7_share_in   ;
assign x0x6x7_share_out         =  x0_share_in & x6_share_in & x7_share_in   ;
assign x1x3x5_share_out         =  x1_share_in & x3_share_in & x5_share_in   ;
assign x1x3x6_share_out         =  x1_share_in & x3_share_in & x6_share_in   ;
assign x1x4x7_share_out         =  x1_share_in & x4_share_in & x7_share_in   ;
assign x2x3x4_share_out         =  x2_share_in & x3_share_in & x4_share_in   ;
assign x2x3x6_share_out         =  x2_share_in & x3_share_in & x6_share_in   ;
assign x3x4x6_share_out         =  x3_share_in & x4_share_in & x6_share_in   ;
assign x3x5x6_share_out         =  x3_share_in & x5_share_in & x6_share_in   ;
assign x0x1x5_share_out         =  x0_share_in & x1_share_in & x5_share_in   ;
assign x0x3x7_share_out         =  x0_share_in & x3_share_in & x7_share_in   ;
assign x1x2x5_share_out         =  x1_share_in & x2_share_in & x5_share_in   ;
assign x1x2x7_share_out         =  x1_share_in & x2_share_in & x7_share_in   ;
assign x1x4x5_share_out         =  x1_share_in & x4_share_in & x5_share_in   ;
assign x1x5x7_share_out         =  x1_share_in & x5_share_in & x7_share_in   ;
assign x2x4x5_share_out         =  x2_share_in & x4_share_in & x5_share_in   ;
assign x3x4x5_share_out         =  x3_share_in & x4_share_in & x5_share_in   ;
assign x4x6x7_share_out         =  x4_share_in & x6_share_in & x7_share_in   ;
assign x1x6x7_share_out         =  x1_share_in & x6_share_in & x7_share_in   ;
assign x4x5x7_share_out         =  x4_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2_share_out         =  x0_share_in & x1_share_in & x2_share_in   ;
assign x0x5x6_share_out         =  x0_share_in & x5_share_in & x6_share_in   ;
assign x2x4x6_share_out         =  x2_share_in & x4_share_in & x6_share_in   ;
assign x0x1x2x3_share_out       =  x0_share_in & x1_share_in & x2_share_in & x3_share_in   ;
assign x0x1x2x5_share_out       =  x0_share_in & x1_share_in & x2_share_in & x5_share_in   ;
assign x0x1x2x6_share_out       =  x0_share_in & x1_share_in & x2_share_in & x6_share_in   ;
assign x0x1x2x7_share_out       =  x0_share_in & x1_share_in & x2_share_in & x7_share_in   ;
assign x0x1x4x5_share_out       =  x0_share_in & x1_share_in & x4_share_in & x5_share_in   ;
assign x0x1x4x7_share_out       =  x0_share_in & x1_share_in & x4_share_in & x7_share_in   ;
assign x0x2x3x5_share_out       =  x0_share_in & x2_share_in & x3_share_in & x5_share_in   ;
assign x0x2x3x7_share_out       =  x0_share_in & x2_share_in & x3_share_in & x7_share_in   ;
assign x0x2x4x5_share_out       =  x0_share_in & x2_share_in & x4_share_in & x5_share_in   ;
assign x0x2x4x7_share_out       =  x0_share_in & x2_share_in & x4_share_in & x7_share_in   ;
assign x0x2x5x6_share_out       =  x0_share_in & x2_share_in & x5_share_in & x6_share_in   ;
assign x0x2x5x7_share_out       =  x0_share_in & x2_share_in & x5_share_in & x7_share_in   ;
assign x0x3x4x6_share_out       =  x0_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x0x3x5x6_share_out       =  x0_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x0x4x5x6_share_out       =  x0_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x4x5x7_share_out       =  x0_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x4x6x7_share_out       =  x0_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x5_share_out       =  x1_share_in & x2_share_in & x3_share_in & x5_share_in   ;
assign x1x2x3x6_share_out       =  x1_share_in & x2_share_in & x3_share_in & x6_share_in   ;
assign x1x2x3x7_share_out       =  x1_share_in & x2_share_in & x3_share_in & x7_share_in   ;
assign x1x2x4x6_share_out       =  x1_share_in & x2_share_in & x4_share_in & x6_share_in   ;
assign x1x2x4x7_share_out       =  x1_share_in & x2_share_in & x4_share_in & x7_share_in   ;
assign x1x2x6x7_share_out       =  x1_share_in & x2_share_in & x6_share_in & x7_share_in   ;
assign x1x3x4x6_share_out       =  x1_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x1x3x6x7_share_out       =  x1_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x1x4x5x6_share_out       =  x1_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x1x4x5x7_share_out       =  x1_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x1x5x6x7_share_out       =  x1_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x2x3x5x7_share_out       =  x2_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x2x3x6x7_share_out       =  x2_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x2x4x5x6_share_out       =  x2_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x2x4x5x7_share_out       =  x2_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x3x5x6x7_share_out       =  x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4_share_out       =  x0_share_in & x1_share_in & x3_share_in & x4_share_in   ;
assign x0x1x3x6_share_out       =  x0_share_in & x1_share_in & x3_share_in & x6_share_in   ;
assign x0x1x5x6_share_out       =  x0_share_in & x1_share_in & x5_share_in & x6_share_in   ;
assign x0x2x3x6_share_out       =  x0_share_in & x2_share_in & x3_share_in & x6_share_in   ;
assign x0x3x4x5_share_out       =  x0_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x1x2x5x6_share_out       =  x1_share_in & x2_share_in & x5_share_in & x6_share_in   ;
assign x1x2x5x7_share_out       =  x1_share_in & x2_share_in & x5_share_in & x7_share_in   ;
assign x1x3x4x5_share_out       =  x1_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x1x3x4x7_share_out       =  x1_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x1x3x5x6_share_out       =  x1_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x1x3x5x7_share_out       =  x1_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x1x4x6x7_share_out       =  x1_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x2x3x4x5_share_out       =  x2_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x2x3x4x7_share_out       =  x2_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x2x4x6x7_share_out       =  x2_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x3x4x5x6_share_out       =  x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x3x4x5x7_share_out       =  x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x3x4x6x7_share_out       =  x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x5_share_out       =  x0_share_in & x1_share_in & x3_share_in & x5_share_in   ;
assign x0x1x4x6_share_out       =  x0_share_in & x1_share_in & x4_share_in & x6_share_in   ;
assign x0x2x3x4_share_out       =  x0_share_in & x2_share_in & x3_share_in & x4_share_in   ;
assign x0x2x4x6_share_out       =  x0_share_in & x2_share_in & x4_share_in & x6_share_in   ;
assign x0x3x4x7_share_out       =  x0_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x3x5x7_share_out       =  x0_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x1x2x3x4_share_out       =  x1_share_in & x2_share_in & x3_share_in & x4_share_in   ;
assign x2x3x4x6_share_out       =  x2_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x2x3x5x6_share_out       =  x2_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x2x5x6x7_share_out       =  x2_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x4x5x6x7_share_out       =  x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x4_share_out       =  x0_share_in & x1_share_in & x2_share_in & x4_share_in   ;
assign x0x1x6x7_share_out       =  x0_share_in & x1_share_in & x6_share_in & x7_share_in   ;
assign x0x2x6x7_share_out       =  x0_share_in & x2_share_in & x6_share_in & x7_share_in   ;
assign x0x3x6x7_share_out       =  x0_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x0x5x6x7_share_out       =  x0_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x4x5_share_out       =  x1_share_in & x2_share_in & x4_share_in & x5_share_in   ;
assign x0x1x3x7_share_out       =  x0_share_in & x1_share_in & x3_share_in & x7_share_in   ;
assign x0x1x5x7_share_out       =  x0_share_in & x1_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2x3x4_share_out     =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in   ;
assign x0x1x2x3x6_share_out     =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x6_share_in   ;
assign x0x1x2x3x7_share_out     =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x7_share_in   ;
assign x0x1x2x4x5_share_out     =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x5_share_in   ;
assign x0x1x2x4x7_share_out     =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x7_share_in   ;
assign x0x1x2x5x7_share_out     =  x0_share_in & x1_share_in & x2_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2x6x7_share_out     =  x0_share_in & x1_share_in & x2_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4x6_share_out     =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x0x1x3x5x6_share_out     =  x0_share_in & x1_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x0x1x3x5x7_share_out     =  x0_share_in & x1_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x0x1x3x6x7_share_out     =  x0_share_in & x1_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x0x1x4x5x6_share_out     =  x0_share_in & x1_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x1x5x6x7_share_out     =  x0_share_in & x1_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x2x3x4x5_share_out     =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x0x2x3x4x6_share_out     =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x0x2x4x5x7_share_out     =  x0_share_in & x2_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x2x4x6x7_share_out     =  x0_share_in & x2_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x3x4x5x6_share_out     =  x0_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x3x4x5x7_share_out     =  x0_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x3x4x6x7_share_out     =  x0_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x3x5x6x7_share_out     =  x0_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x5x6_share_out     =  x1_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x1x2x3x5x7_share_out     =  x1_share_in & x2_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x1x2x4x5x6_share_out     =  x1_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x1x2x4x6x7_share_out     =  x1_share_in & x2_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x5x6x7_share_out     =  x1_share_in & x2_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x3x4x5x7_share_out     =  x1_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x2x3x4x5x6_share_out     =  x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x2x3x4x5x7_share_out     =  x2_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x2x4x5x6x7_share_out     =  x2_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x4x6_share_out     =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x6_share_in   ;
assign x0x1x3x4x7_share_out     =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x2x3x4x7_share_out     =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x2x3x5x7_share_out     =  x0_share_in & x2_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x0x2x3x6x7_share_out     =  x0_share_in & x2_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x0x2x4x5x6_share_out     =  x0_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x2x5x6x7_share_out     =  x0_share_in & x2_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x4x5x6x7_share_out     =  x0_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x6_share_out     =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x1x3x4x5x6_share_out     =  x1_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x2x3x4x6x7_share_out     =  x2_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x5_share_out     =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x5_share_in   ;
assign x0x1x4x6x7_share_out     =  x0_share_in & x1_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x5_share_out     =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x1x2x3x6x7_share_out     =  x1_share_in & x2_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x1x2x4x5x7_share_out     =  x1_share_in & x2_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x1x3x4x6x7_share_out     =  x1_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x3x5x6x7_share_out     =  x1_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x4x5x6x7_share_out     =  x1_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x2x3x5x6x7_share_out     =  x2_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x3x4x5x6x7_share_out     =  x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x5x6_share_out     =  x0_share_in & x1_share_in & x2_share_in & x5_share_in & x6_share_in   ;
assign x0x1x3x4x5_share_out     =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x0x1x4x5x7_share_out     =  x0_share_in & x1_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x2x3x5x6_share_out     =  x0_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x1x2x3x4x7_share_out     =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x1x2x3x4x6_share_out   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x0x1x2x3x4x7_share_out   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x1x2x3x5x7_share_out   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2x3x6x7_share_out   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x4x5x7_share_out   =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2x5x6x7_share_out   =  x0_share_in & x1_share_in & x2_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4x6x7_share_out   =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x4x5x6x7_share_out   =  x0_share_in & x1_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x2x3x4x5x6_share_out   =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x2x3x4x5x7_share_out   =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x2x3x5x6x7_share_out   =  x0_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x6x7_share_out   =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x4x5x6x7_share_out   =  x1_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x3x4x5x6x7_share_out   =  x1_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x2x3x4x5x6x7_share_out   =  x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x5x6_share_out   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x0x1x2x4x6x7_share_out   =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4x5x6_share_out   =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x2x3x4x6x7_share_out   =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x5x6_share_out   =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x1x2x3x5x6x7_share_out   =  x1_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x4x5_share_out   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x0x1x2x4x5x6_share_out   =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x1x3x4x5x7_share_out   =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x1x3x5x6x7_share_out   =  x0_share_in & x1_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x2x4x5x6x7_share_out   =  x0_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x5x7_share_out   =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x3x4x5x6x7_share_out   =  x0_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x4x6x7_share_out =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x4x5x6x7_share_out =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x2x3x4x5x6x7_share_out =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x5x6x7_share_out =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4x5x6x7_share_out =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x5x6x7_share_out =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x4x5x6_share_out =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x1x2x3x4x5x7_share_out =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;

endmodule