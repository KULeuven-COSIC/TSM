`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 02/22/2025
// Design Name: Second-Order Masked AES S-Box
// Module Name: AES_sbox_secondorder_threeregstages
// Description: Implements a second-order masked AES S-Box using HO-TSM2 with three register stages.
// Dependencies: None
// Revision: 0.01 - Initial version
//////////////////////////////////////////////////////////////////////////////////

module AES_sbox_secondorder_threeregstages ( clk, 
rand_bit_cycle1, rand_bit_cycle2, rand_bit_cycle3, 
sbox_input_share1, sbox_input_share2, sbox_input_share3,
output_sbox_share1, output_sbox_share2, output_sbox_share3
);


input clk;
input [54:1] rand_bit_cycle1;
input [60:1] rand_bit_cycle2;
input [24:1] rand_bit_cycle3;

input [7:0] sbox_input_share1, sbox_input_share2, sbox_input_share3;
output [7:0] output_sbox_share1, output_sbox_share2, output_sbox_share3;


wire x0_input_share1 = sbox_input_share1[0];
wire x1_input_share1 = sbox_input_share1[1];
wire x2_input_share1 = sbox_input_share1[2];
wire x3_input_share1 = sbox_input_share1[3];
wire x4_input_share1 = sbox_input_share1[4];
wire x5_input_share1 = sbox_input_share1[5];
wire x6_input_share1 = sbox_input_share1[6];
wire x7_input_share1 = sbox_input_share1[7];

wire x0_input_share2 = sbox_input_share2[0];
wire x1_input_share2 = sbox_input_share2[1];
wire x2_input_share2 = sbox_input_share2[2];
wire x3_input_share2 = sbox_input_share2[3];
wire x4_input_share2 = sbox_input_share2[4];
wire x5_input_share2 = sbox_input_share2[5];
wire x6_input_share2 = sbox_input_share2[6];
wire x7_input_share2 = sbox_input_share2[7];

wire x0_input_share3 = sbox_input_share3[0];
wire x1_input_share3 = sbox_input_share3[1];
wire x2_input_share3 = sbox_input_share3[2];
wire x3_input_share3 = sbox_input_share3[3];
wire x4_input_share3 = sbox_input_share3[4];
wire x5_input_share3 = sbox_input_share3[5];
wire x6_input_share3 = sbox_input_share3[6];
wire x7_input_share3 = sbox_input_share3[7];


HO_TSM2_fourinput_secondorder_block first_module(clk, rand_bit_cycle1[27:1] , rand_bit_cycle2[30:1]  , x0_input_share1, x1_input_share1, x2_input_share1, x3_input_share1,  x0_input_share2, x1_input_share2, x2_input_share2, x3_input_share2,  x0_input_share3, x1_input_share3, x2_input_share3, x3_input_share3, output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 , output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 , output_x0_share3, output_x1_share3, output_x2_share3, output_x3_share3, output_x0x1_share3, output_x0x2_share3, output_x0x3_share3, output_x1x2_share3, output_x1x3_share3, output_x2x3_share3, output_x0x1x2_share3, output_x0x1x3_share3, output_x0x2x3_share3, output_x1x2x3_share3, output_x0x1x2x3_share3 );
HO_TSM2_fourinput_secondorder_block secon_module(clk, rand_bit_cycle1[54:28], rand_bit_cycle2[60:31] , x4_input_share1, x5_input_share1, x6_input_share1, x7_input_share1,  x4_input_share2, x5_input_share2, x6_input_share2, x7_input_share2,  x4_input_share3, x5_input_share3, x6_input_share3, x7_input_share3, output_x4_share1, output_x5_share1, output_x6_share1, output_x7_share1, output_x4x5_share1, output_x4x6_share1, output_x4x7_share1, output_x5x6_share1, output_x5x7_share1, output_x6x7_share1, output_x4x5x6_share1, output_x4x5x7_share1, output_x4x6x7_share1, output_x5x6x7_share1, output_x4x5x6x7_share1 , output_x4_share2, output_x5_share2, output_x6_share2, output_x7_share2, output_x4x5_share2, output_x4x6_share2, output_x4x7_share2, output_x5x6_share2, output_x5x7_share2, output_x6x7_share2, output_x4x5x6_share2, output_x4x5x7_share2, output_x4x6x7_share2, output_x5x6x7_share2, output_x4x5x6x7_share2 , output_x4_share3, output_x5_share3, output_x6_share3, output_x7_share3, output_x4x5_share3, output_x4x6_share3, output_x4x7_share3, output_x5x6_share3, output_x5x7_share3, output_x6x7_share3, output_x4x5x6_share3, output_x4x5x7_share3, output_x4x6x7_share3, output_x5x6x7_share3, output_x4x5x6x7_share3 );


wire [24:1] rand_bit_second;
assign rand_bit_second = rand_bit_cycle3;



wire output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1 ;

wire output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2 ;

wire output_sum_secondmodule_equation_num_0_index_0_share3, output_sum_secondmodule_equation_num_0_index_1_share3, output_sum_secondmodule_equation_num_0_index_2_share3, output_sum_secondmodule_equation_num_0_index_3_share3, output_sum_secondmodule_equation_num_0_index_4_share3, output_sum_secondmodule_equation_num_0_index_5_share3, output_sum_secondmodule_equation_num_0_index_6_share3, output_sum_secondmodule_equation_num_0_index_7_share3, output_sum_secondmodule_equation_num_0_index_8_share3, output_sum_secondmodule_equation_num_0_index_9_share3, output_sum_secondmodule_equation_num_0_index_10_share3, output_sum_secondmodule_equation_num_0_index_11_share3, output_sum_secondmodule_equation_num_0_index_12_share3, output_sum_secondmodule_equation_num_0_index_13_share3, output_sum_secondmodule_equation_num_0_index_14_share3,
output_sum_secondmodule_equation_num_1_index_0_share3, output_sum_secondmodule_equation_num_1_index_1_share3, output_sum_secondmodule_equation_num_1_index_2_share3, output_sum_secondmodule_equation_num_1_index_3_share3, output_sum_secondmodule_equation_num_1_index_4_share3, output_sum_secondmodule_equation_num_1_index_5_share3, output_sum_secondmodule_equation_num_1_index_6_share3, output_sum_secondmodule_equation_num_1_index_7_share3, output_sum_secondmodule_equation_num_1_index_8_share3, output_sum_secondmodule_equation_num_1_index_9_share3, output_sum_secondmodule_equation_num_1_index_10_share3, output_sum_secondmodule_equation_num_1_index_11_share3, output_sum_secondmodule_equation_num_1_index_12_share3, output_sum_secondmodule_equation_num_1_index_13_share3, output_sum_secondmodule_equation_num_1_index_14_share3,
output_sum_secondmodule_equation_num_2_index_0_share3, output_sum_secondmodule_equation_num_2_index_1_share3, output_sum_secondmodule_equation_num_2_index_2_share3, output_sum_secondmodule_equation_num_2_index_3_share3, output_sum_secondmodule_equation_num_2_index_4_share3, output_sum_secondmodule_equation_num_2_index_5_share3, output_sum_secondmodule_equation_num_2_index_6_share3, output_sum_secondmodule_equation_num_2_index_7_share3, output_sum_secondmodule_equation_num_2_index_8_share3, output_sum_secondmodule_equation_num_2_index_9_share3, output_sum_secondmodule_equation_num_2_index_10_share3, output_sum_secondmodule_equation_num_2_index_11_share3, output_sum_secondmodule_equation_num_2_index_12_share3, output_sum_secondmodule_equation_num_2_index_13_share3, output_sum_secondmodule_equation_num_2_index_14_share3,
output_sum_secondmodule_equation_num_3_index_0_share3, output_sum_secondmodule_equation_num_3_index_1_share3, output_sum_secondmodule_equation_num_3_index_2_share3, output_sum_secondmodule_equation_num_3_index_3_share3, output_sum_secondmodule_equation_num_3_index_4_share3, output_sum_secondmodule_equation_num_3_index_5_share3, output_sum_secondmodule_equation_num_3_index_6_share3, output_sum_secondmodule_equation_num_3_index_7_share3, output_sum_secondmodule_equation_num_3_index_8_share3, output_sum_secondmodule_equation_num_3_index_9_share3, output_sum_secondmodule_equation_num_3_index_10_share3, output_sum_secondmodule_equation_num_3_index_11_share3, output_sum_secondmodule_equation_num_3_index_12_share3, output_sum_secondmodule_equation_num_3_index_13_share3, output_sum_secondmodule_equation_num_3_index_14_share3,
output_sum_secondmodule_equation_num_4_index_0_share3, output_sum_secondmodule_equation_num_4_index_1_share3, output_sum_secondmodule_equation_num_4_index_2_share3, output_sum_secondmodule_equation_num_4_index_3_share3, output_sum_secondmodule_equation_num_4_index_4_share3, output_sum_secondmodule_equation_num_4_index_5_share3, output_sum_secondmodule_equation_num_4_index_6_share3, output_sum_secondmodule_equation_num_4_index_7_share3, output_sum_secondmodule_equation_num_4_index_8_share3, output_sum_secondmodule_equation_num_4_index_9_share3, output_sum_secondmodule_equation_num_4_index_10_share3, output_sum_secondmodule_equation_num_4_index_11_share3, output_sum_secondmodule_equation_num_4_index_12_share3, output_sum_secondmodule_equation_num_4_index_13_share3, output_sum_secondmodule_equation_num_4_index_14_share3,
output_sum_secondmodule_equation_num_5_index_0_share3, output_sum_secondmodule_equation_num_5_index_1_share3, output_sum_secondmodule_equation_num_5_index_2_share3, output_sum_secondmodule_equation_num_5_index_3_share3, output_sum_secondmodule_equation_num_5_index_4_share3, output_sum_secondmodule_equation_num_5_index_5_share3, output_sum_secondmodule_equation_num_5_index_6_share3, output_sum_secondmodule_equation_num_5_index_7_share3, output_sum_secondmodule_equation_num_5_index_8_share3, output_sum_secondmodule_equation_num_5_index_9_share3, output_sum_secondmodule_equation_num_5_index_10_share3, output_sum_secondmodule_equation_num_5_index_11_share3, output_sum_secondmodule_equation_num_5_index_12_share3, output_sum_secondmodule_equation_num_5_index_13_share3, output_sum_secondmodule_equation_num_5_index_14_share3,
output_sum_secondmodule_equation_num_6_index_0_share3, output_sum_secondmodule_equation_num_6_index_1_share3, output_sum_secondmodule_equation_num_6_index_2_share3, output_sum_secondmodule_equation_num_6_index_3_share3, output_sum_secondmodule_equation_num_6_index_4_share3, output_sum_secondmodule_equation_num_6_index_5_share3, output_sum_secondmodule_equation_num_6_index_6_share3, output_sum_secondmodule_equation_num_6_index_7_share3, output_sum_secondmodule_equation_num_6_index_8_share3, output_sum_secondmodule_equation_num_6_index_9_share3, output_sum_secondmodule_equation_num_6_index_10_share3, output_sum_secondmodule_equation_num_6_index_11_share3, output_sum_secondmodule_equation_num_6_index_12_share3, output_sum_secondmodule_equation_num_6_index_13_share3, output_sum_secondmodule_equation_num_6_index_14_share3,
output_sum_secondmodule_equation_num_7_index_0_share3, output_sum_secondmodule_equation_num_7_index_1_share3, output_sum_secondmodule_equation_num_7_index_2_share3, output_sum_secondmodule_equation_num_7_index_3_share3, output_sum_secondmodule_equation_num_7_index_4_share3, output_sum_secondmodule_equation_num_7_index_5_share3, output_sum_secondmodule_equation_num_7_index_6_share3, output_sum_secondmodule_equation_num_7_index_7_share3, output_sum_secondmodule_equation_num_7_index_8_share3, output_sum_secondmodule_equation_num_7_index_9_share3, output_sum_secondmodule_equation_num_7_index_10_share3, output_sum_secondmodule_equation_num_7_index_11_share3, output_sum_secondmodule_equation_num_7_index_12_share3, output_sum_secondmodule_equation_num_7_index_13_share3, output_sum_secondmodule_equation_num_7_index_14_share3 ;

sum_of_second_module_outputs instance_share1 (
    output_x4_share1 ,  output_x5_share1 ,  output_x6_share1 ,  output_x7_share1 ,  output_x4x5_share1 ,  output_x4x6_share1 ,  output_x4x7_share1 ,  output_x5x6_share1 ,  output_x5x7_share1 ,  output_x6x7_share1 ,  output_x4x5x6_share1 ,  output_x4x5x7_share1 ,  output_x4x6x7_share1 ,  output_x5x6x7_share1 ,  output_x4x5x6x7_share1,
output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1

);

sum_of_second_module_outputs instance_share2 (
    output_x4_share2 ,  output_x5_share2 ,  output_x6_share2 ,  output_x7_share2 ,  output_x4x5_share2 ,  output_x4x6_share2 ,  output_x4x7_share2 ,  output_x5x6_share2 ,  output_x5x7_share2 ,  output_x6x7_share2 ,  output_x4x5x6_share2 ,  output_x4x5x7_share2 ,  output_x4x6x7_share2 ,  output_x5x6x7_share2 ,  output_x4x5x6x7_share2,
output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2

);

sum_of_second_module_outputs instance_share3 (
    output_x4_share3 ,  output_x5_share3 ,  output_x6_share3 ,  output_x7_share3 ,  output_x4x5_share3 ,  output_x4x6_share3 ,  output_x4x7_share3 ,  output_x5x6_share3 ,  output_x5x7_share3 ,  output_x6x7_share3 ,  output_x4x5x6_share3 ,  output_x4x5x7_share3 ,  output_x4x6x7_share3 ,  output_x5x6x7_share3 ,  output_x4x5x6x7_share3,
output_sum_secondmodule_equation_num_0_index_0_share3, output_sum_secondmodule_equation_num_0_index_1_share3, output_sum_secondmodule_equation_num_0_index_2_share3, output_sum_secondmodule_equation_num_0_index_3_share3, output_sum_secondmodule_equation_num_0_index_4_share3, output_sum_secondmodule_equation_num_0_index_5_share3, output_sum_secondmodule_equation_num_0_index_6_share3, output_sum_secondmodule_equation_num_0_index_7_share3, output_sum_secondmodule_equation_num_0_index_8_share3, output_sum_secondmodule_equation_num_0_index_9_share3, output_sum_secondmodule_equation_num_0_index_10_share3, output_sum_secondmodule_equation_num_0_index_11_share3, output_sum_secondmodule_equation_num_0_index_12_share3, output_sum_secondmodule_equation_num_0_index_13_share3, output_sum_secondmodule_equation_num_0_index_14_share3,
output_sum_secondmodule_equation_num_1_index_0_share3, output_sum_secondmodule_equation_num_1_index_1_share3, output_sum_secondmodule_equation_num_1_index_2_share3, output_sum_secondmodule_equation_num_1_index_3_share3, output_sum_secondmodule_equation_num_1_index_4_share3, output_sum_secondmodule_equation_num_1_index_5_share3, output_sum_secondmodule_equation_num_1_index_6_share3, output_sum_secondmodule_equation_num_1_index_7_share3, output_sum_secondmodule_equation_num_1_index_8_share3, output_sum_secondmodule_equation_num_1_index_9_share3, output_sum_secondmodule_equation_num_1_index_10_share3, output_sum_secondmodule_equation_num_1_index_11_share3, output_sum_secondmodule_equation_num_1_index_12_share3, output_sum_secondmodule_equation_num_1_index_13_share3, output_sum_secondmodule_equation_num_1_index_14_share3,
output_sum_secondmodule_equation_num_2_index_0_share3, output_sum_secondmodule_equation_num_2_index_1_share3, output_sum_secondmodule_equation_num_2_index_2_share3, output_sum_secondmodule_equation_num_2_index_3_share3, output_sum_secondmodule_equation_num_2_index_4_share3, output_sum_secondmodule_equation_num_2_index_5_share3, output_sum_secondmodule_equation_num_2_index_6_share3, output_sum_secondmodule_equation_num_2_index_7_share3, output_sum_secondmodule_equation_num_2_index_8_share3, output_sum_secondmodule_equation_num_2_index_9_share3, output_sum_secondmodule_equation_num_2_index_10_share3, output_sum_secondmodule_equation_num_2_index_11_share3, output_sum_secondmodule_equation_num_2_index_12_share3, output_sum_secondmodule_equation_num_2_index_13_share3, output_sum_secondmodule_equation_num_2_index_14_share3,
output_sum_secondmodule_equation_num_3_index_0_share3, output_sum_secondmodule_equation_num_3_index_1_share3, output_sum_secondmodule_equation_num_3_index_2_share3, output_sum_secondmodule_equation_num_3_index_3_share3, output_sum_secondmodule_equation_num_3_index_4_share3, output_sum_secondmodule_equation_num_3_index_5_share3, output_sum_secondmodule_equation_num_3_index_6_share3, output_sum_secondmodule_equation_num_3_index_7_share3, output_sum_secondmodule_equation_num_3_index_8_share3, output_sum_secondmodule_equation_num_3_index_9_share3, output_sum_secondmodule_equation_num_3_index_10_share3, output_sum_secondmodule_equation_num_3_index_11_share3, output_sum_secondmodule_equation_num_3_index_12_share3, output_sum_secondmodule_equation_num_3_index_13_share3, output_sum_secondmodule_equation_num_3_index_14_share3,
output_sum_secondmodule_equation_num_4_index_0_share3, output_sum_secondmodule_equation_num_4_index_1_share3, output_sum_secondmodule_equation_num_4_index_2_share3, output_sum_secondmodule_equation_num_4_index_3_share3, output_sum_secondmodule_equation_num_4_index_4_share3, output_sum_secondmodule_equation_num_4_index_5_share3, output_sum_secondmodule_equation_num_4_index_6_share3, output_sum_secondmodule_equation_num_4_index_7_share3, output_sum_secondmodule_equation_num_4_index_8_share3, output_sum_secondmodule_equation_num_4_index_9_share3, output_sum_secondmodule_equation_num_4_index_10_share3, output_sum_secondmodule_equation_num_4_index_11_share3, output_sum_secondmodule_equation_num_4_index_12_share3, output_sum_secondmodule_equation_num_4_index_13_share3, output_sum_secondmodule_equation_num_4_index_14_share3,
output_sum_secondmodule_equation_num_5_index_0_share3, output_sum_secondmodule_equation_num_5_index_1_share3, output_sum_secondmodule_equation_num_5_index_2_share3, output_sum_secondmodule_equation_num_5_index_3_share3, output_sum_secondmodule_equation_num_5_index_4_share3, output_sum_secondmodule_equation_num_5_index_5_share3, output_sum_secondmodule_equation_num_5_index_6_share3, output_sum_secondmodule_equation_num_5_index_7_share3, output_sum_secondmodule_equation_num_5_index_8_share3, output_sum_secondmodule_equation_num_5_index_9_share3, output_sum_secondmodule_equation_num_5_index_10_share3, output_sum_secondmodule_equation_num_5_index_11_share3, output_sum_secondmodule_equation_num_5_index_12_share3, output_sum_secondmodule_equation_num_5_index_13_share3, output_sum_secondmodule_equation_num_5_index_14_share3,
output_sum_secondmodule_equation_num_6_index_0_share3, output_sum_secondmodule_equation_num_6_index_1_share3, output_sum_secondmodule_equation_num_6_index_2_share3, output_sum_secondmodule_equation_num_6_index_3_share3, output_sum_secondmodule_equation_num_6_index_4_share3, output_sum_secondmodule_equation_num_6_index_5_share3, output_sum_secondmodule_equation_num_6_index_6_share3, output_sum_secondmodule_equation_num_6_index_7_share3, output_sum_secondmodule_equation_num_6_index_8_share3, output_sum_secondmodule_equation_num_6_index_9_share3, output_sum_secondmodule_equation_num_6_index_10_share3, output_sum_secondmodule_equation_num_6_index_11_share3, output_sum_secondmodule_equation_num_6_index_12_share3, output_sum_secondmodule_equation_num_6_index_13_share3, output_sum_secondmodule_equation_num_6_index_14_share3,
output_sum_secondmodule_equation_num_7_index_0_share3, output_sum_secondmodule_equation_num_7_index_1_share3, output_sum_secondmodule_equation_num_7_index_2_share3, output_sum_secondmodule_equation_num_7_index_3_share3, output_sum_secondmodule_equation_num_7_index_4_share3, output_sum_secondmodule_equation_num_7_index_5_share3, output_sum_secondmodule_equation_num_7_index_6_share3, output_sum_secondmodule_equation_num_7_index_7_share3, output_sum_secondmodule_equation_num_7_index_8_share3, output_sum_secondmodule_equation_num_7_index_9_share3, output_sum_secondmodule_equation_num_7_index_10_share3, output_sum_secondmodule_equation_num_7_index_11_share3, output_sum_secondmodule_equation_num_7_index_12_share3, output_sum_secondmodule_equation_num_7_index_13_share3, output_sum_secondmodule_equation_num_7_index_14_share3

);

// DOM-indep multiplications, cross module terms


cross_module_multiplication inst_domain_1 (
output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 , 
output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1,
cross_module_equation_num0_domain_1, cross_module_equation_num1_domain_1, cross_module_equation_num2_domain_1, cross_module_equation_num3_domain_1,cross_module_equation_num4_domain_1,cross_module_equation_num5_domain_1,cross_module_equation_num6_domain_1,cross_module_equation_num7_domain_1
);


cross_module_multiplication inst_domain_2 (
output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 , 
output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2,
cross_module_equation_num0_domain_2, cross_module_equation_num1_domain_2, cross_module_equation_num2_domain_2, cross_module_equation_num3_domain_2,cross_module_equation_num4_domain_2,cross_module_equation_num5_domain_2,cross_module_equation_num6_domain_2,cross_module_equation_num7_domain_2
);


cross_module_multiplication inst_domain_3 (
output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 , 
output_sum_secondmodule_equation_num_0_index_0_share3, output_sum_secondmodule_equation_num_0_index_1_share3, output_sum_secondmodule_equation_num_0_index_2_share3, output_sum_secondmodule_equation_num_0_index_3_share3, output_sum_secondmodule_equation_num_0_index_4_share3, output_sum_secondmodule_equation_num_0_index_5_share3, output_sum_secondmodule_equation_num_0_index_6_share3, output_sum_secondmodule_equation_num_0_index_7_share3, output_sum_secondmodule_equation_num_0_index_8_share3, output_sum_secondmodule_equation_num_0_index_9_share3, output_sum_secondmodule_equation_num_0_index_10_share3, output_sum_secondmodule_equation_num_0_index_11_share3, output_sum_secondmodule_equation_num_0_index_12_share3, output_sum_secondmodule_equation_num_0_index_13_share3, output_sum_secondmodule_equation_num_0_index_14_share3,
output_sum_secondmodule_equation_num_1_index_0_share3, output_sum_secondmodule_equation_num_1_index_1_share3, output_sum_secondmodule_equation_num_1_index_2_share3, output_sum_secondmodule_equation_num_1_index_3_share3, output_sum_secondmodule_equation_num_1_index_4_share3, output_sum_secondmodule_equation_num_1_index_5_share3, output_sum_secondmodule_equation_num_1_index_6_share3, output_sum_secondmodule_equation_num_1_index_7_share3, output_sum_secondmodule_equation_num_1_index_8_share3, output_sum_secondmodule_equation_num_1_index_9_share3, output_sum_secondmodule_equation_num_1_index_10_share3, output_sum_secondmodule_equation_num_1_index_11_share3, output_sum_secondmodule_equation_num_1_index_12_share3, output_sum_secondmodule_equation_num_1_index_13_share3, output_sum_secondmodule_equation_num_1_index_14_share3,
output_sum_secondmodule_equation_num_2_index_0_share3, output_sum_secondmodule_equation_num_2_index_1_share3, output_sum_secondmodule_equation_num_2_index_2_share3, output_sum_secondmodule_equation_num_2_index_3_share3, output_sum_secondmodule_equation_num_2_index_4_share3, output_sum_secondmodule_equation_num_2_index_5_share3, output_sum_secondmodule_equation_num_2_index_6_share3, output_sum_secondmodule_equation_num_2_index_7_share3, output_sum_secondmodule_equation_num_2_index_8_share3, output_sum_secondmodule_equation_num_2_index_9_share3, output_sum_secondmodule_equation_num_2_index_10_share3, output_sum_secondmodule_equation_num_2_index_11_share3, output_sum_secondmodule_equation_num_2_index_12_share3, output_sum_secondmodule_equation_num_2_index_13_share3, output_sum_secondmodule_equation_num_2_index_14_share3,
output_sum_secondmodule_equation_num_3_index_0_share3, output_sum_secondmodule_equation_num_3_index_1_share3, output_sum_secondmodule_equation_num_3_index_2_share3, output_sum_secondmodule_equation_num_3_index_3_share3, output_sum_secondmodule_equation_num_3_index_4_share3, output_sum_secondmodule_equation_num_3_index_5_share3, output_sum_secondmodule_equation_num_3_index_6_share3, output_sum_secondmodule_equation_num_3_index_7_share3, output_sum_secondmodule_equation_num_3_index_8_share3, output_sum_secondmodule_equation_num_3_index_9_share3, output_sum_secondmodule_equation_num_3_index_10_share3, output_sum_secondmodule_equation_num_3_index_11_share3, output_sum_secondmodule_equation_num_3_index_12_share3, output_sum_secondmodule_equation_num_3_index_13_share3, output_sum_secondmodule_equation_num_3_index_14_share3,
output_sum_secondmodule_equation_num_4_index_0_share3, output_sum_secondmodule_equation_num_4_index_1_share3, output_sum_secondmodule_equation_num_4_index_2_share3, output_sum_secondmodule_equation_num_4_index_3_share3, output_sum_secondmodule_equation_num_4_index_4_share3, output_sum_secondmodule_equation_num_4_index_5_share3, output_sum_secondmodule_equation_num_4_index_6_share3, output_sum_secondmodule_equation_num_4_index_7_share3, output_sum_secondmodule_equation_num_4_index_8_share3, output_sum_secondmodule_equation_num_4_index_9_share3, output_sum_secondmodule_equation_num_4_index_10_share3, output_sum_secondmodule_equation_num_4_index_11_share3, output_sum_secondmodule_equation_num_4_index_12_share3, output_sum_secondmodule_equation_num_4_index_13_share3, output_sum_secondmodule_equation_num_4_index_14_share3,
output_sum_secondmodule_equation_num_5_index_0_share3, output_sum_secondmodule_equation_num_5_index_1_share3, output_sum_secondmodule_equation_num_5_index_2_share3, output_sum_secondmodule_equation_num_5_index_3_share3, output_sum_secondmodule_equation_num_5_index_4_share3, output_sum_secondmodule_equation_num_5_index_5_share3, output_sum_secondmodule_equation_num_5_index_6_share3, output_sum_secondmodule_equation_num_5_index_7_share3, output_sum_secondmodule_equation_num_5_index_8_share3, output_sum_secondmodule_equation_num_5_index_9_share3, output_sum_secondmodule_equation_num_5_index_10_share3, output_sum_secondmodule_equation_num_5_index_11_share3, output_sum_secondmodule_equation_num_5_index_12_share3, output_sum_secondmodule_equation_num_5_index_13_share3, output_sum_secondmodule_equation_num_5_index_14_share3,
output_sum_secondmodule_equation_num_6_index_0_share3, output_sum_secondmodule_equation_num_6_index_1_share3, output_sum_secondmodule_equation_num_6_index_2_share3, output_sum_secondmodule_equation_num_6_index_3_share3, output_sum_secondmodule_equation_num_6_index_4_share3, output_sum_secondmodule_equation_num_6_index_5_share3, output_sum_secondmodule_equation_num_6_index_6_share3, output_sum_secondmodule_equation_num_6_index_7_share3, output_sum_secondmodule_equation_num_6_index_8_share3, output_sum_secondmodule_equation_num_6_index_9_share3, output_sum_secondmodule_equation_num_6_index_10_share3, output_sum_secondmodule_equation_num_6_index_11_share3, output_sum_secondmodule_equation_num_6_index_12_share3, output_sum_secondmodule_equation_num_6_index_13_share3, output_sum_secondmodule_equation_num_6_index_14_share3,
output_sum_secondmodule_equation_num_7_index_0_share3, output_sum_secondmodule_equation_num_7_index_1_share3, output_sum_secondmodule_equation_num_7_index_2_share3, output_sum_secondmodule_equation_num_7_index_3_share3, output_sum_secondmodule_equation_num_7_index_4_share3, output_sum_secondmodule_equation_num_7_index_5_share3, output_sum_secondmodule_equation_num_7_index_6_share3, output_sum_secondmodule_equation_num_7_index_7_share3, output_sum_secondmodule_equation_num_7_index_8_share3, output_sum_secondmodule_equation_num_7_index_9_share3, output_sum_secondmodule_equation_num_7_index_10_share3, output_sum_secondmodule_equation_num_7_index_11_share3, output_sum_secondmodule_equation_num_7_index_12_share3, output_sum_secondmodule_equation_num_7_index_13_share3, output_sum_secondmodule_equation_num_7_index_14_share3,
cross_module_equation_num0_domain_3, cross_module_equation_num1_domain_3, cross_module_equation_num2_domain_3, cross_module_equation_num3_domain_3,cross_module_equation_num4_domain_3,cross_module_equation_num5_domain_3,cross_module_equation_num6_domain_3,cross_module_equation_num7_domain_3
);


cross_module_multiplication inst_domain_4 (
output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 , 
output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1,
cross_module_equation_num0_domain_4, cross_module_equation_num1_domain_4, cross_module_equation_num2_domain_4, cross_module_equation_num3_domain_4,cross_module_equation_num4_domain_4,cross_module_equation_num5_domain_4,cross_module_equation_num6_domain_4,cross_module_equation_num7_domain_4
);


cross_module_multiplication inst_domain_5 (
output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 , 
output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2,
cross_module_equation_num0_domain_5, cross_module_equation_num1_domain_5, cross_module_equation_num2_domain_5, cross_module_equation_num3_domain_5,cross_module_equation_num4_domain_5,cross_module_equation_num5_domain_5,cross_module_equation_num6_domain_5,cross_module_equation_num7_domain_5
);


cross_module_multiplication inst_domain_6 (
output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 , 
output_sum_secondmodule_equation_num_0_index_0_share3, output_sum_secondmodule_equation_num_0_index_1_share3, output_sum_secondmodule_equation_num_0_index_2_share3, output_sum_secondmodule_equation_num_0_index_3_share3, output_sum_secondmodule_equation_num_0_index_4_share3, output_sum_secondmodule_equation_num_0_index_5_share3, output_sum_secondmodule_equation_num_0_index_6_share3, output_sum_secondmodule_equation_num_0_index_7_share3, output_sum_secondmodule_equation_num_0_index_8_share3, output_sum_secondmodule_equation_num_0_index_9_share3, output_sum_secondmodule_equation_num_0_index_10_share3, output_sum_secondmodule_equation_num_0_index_11_share3, output_sum_secondmodule_equation_num_0_index_12_share3, output_sum_secondmodule_equation_num_0_index_13_share3, output_sum_secondmodule_equation_num_0_index_14_share3,
output_sum_secondmodule_equation_num_1_index_0_share3, output_sum_secondmodule_equation_num_1_index_1_share3, output_sum_secondmodule_equation_num_1_index_2_share3, output_sum_secondmodule_equation_num_1_index_3_share3, output_sum_secondmodule_equation_num_1_index_4_share3, output_sum_secondmodule_equation_num_1_index_5_share3, output_sum_secondmodule_equation_num_1_index_6_share3, output_sum_secondmodule_equation_num_1_index_7_share3, output_sum_secondmodule_equation_num_1_index_8_share3, output_sum_secondmodule_equation_num_1_index_9_share3, output_sum_secondmodule_equation_num_1_index_10_share3, output_sum_secondmodule_equation_num_1_index_11_share3, output_sum_secondmodule_equation_num_1_index_12_share3, output_sum_secondmodule_equation_num_1_index_13_share3, output_sum_secondmodule_equation_num_1_index_14_share3,
output_sum_secondmodule_equation_num_2_index_0_share3, output_sum_secondmodule_equation_num_2_index_1_share3, output_sum_secondmodule_equation_num_2_index_2_share3, output_sum_secondmodule_equation_num_2_index_3_share3, output_sum_secondmodule_equation_num_2_index_4_share3, output_sum_secondmodule_equation_num_2_index_5_share3, output_sum_secondmodule_equation_num_2_index_6_share3, output_sum_secondmodule_equation_num_2_index_7_share3, output_sum_secondmodule_equation_num_2_index_8_share3, output_sum_secondmodule_equation_num_2_index_9_share3, output_sum_secondmodule_equation_num_2_index_10_share3, output_sum_secondmodule_equation_num_2_index_11_share3, output_sum_secondmodule_equation_num_2_index_12_share3, output_sum_secondmodule_equation_num_2_index_13_share3, output_sum_secondmodule_equation_num_2_index_14_share3,
output_sum_secondmodule_equation_num_3_index_0_share3, output_sum_secondmodule_equation_num_3_index_1_share3, output_sum_secondmodule_equation_num_3_index_2_share3, output_sum_secondmodule_equation_num_3_index_3_share3, output_sum_secondmodule_equation_num_3_index_4_share3, output_sum_secondmodule_equation_num_3_index_5_share3, output_sum_secondmodule_equation_num_3_index_6_share3, output_sum_secondmodule_equation_num_3_index_7_share3, output_sum_secondmodule_equation_num_3_index_8_share3, output_sum_secondmodule_equation_num_3_index_9_share3, output_sum_secondmodule_equation_num_3_index_10_share3, output_sum_secondmodule_equation_num_3_index_11_share3, output_sum_secondmodule_equation_num_3_index_12_share3, output_sum_secondmodule_equation_num_3_index_13_share3, output_sum_secondmodule_equation_num_3_index_14_share3,
output_sum_secondmodule_equation_num_4_index_0_share3, output_sum_secondmodule_equation_num_4_index_1_share3, output_sum_secondmodule_equation_num_4_index_2_share3, output_sum_secondmodule_equation_num_4_index_3_share3, output_sum_secondmodule_equation_num_4_index_4_share3, output_sum_secondmodule_equation_num_4_index_5_share3, output_sum_secondmodule_equation_num_4_index_6_share3, output_sum_secondmodule_equation_num_4_index_7_share3, output_sum_secondmodule_equation_num_4_index_8_share3, output_sum_secondmodule_equation_num_4_index_9_share3, output_sum_secondmodule_equation_num_4_index_10_share3, output_sum_secondmodule_equation_num_4_index_11_share3, output_sum_secondmodule_equation_num_4_index_12_share3, output_sum_secondmodule_equation_num_4_index_13_share3, output_sum_secondmodule_equation_num_4_index_14_share3,
output_sum_secondmodule_equation_num_5_index_0_share3, output_sum_secondmodule_equation_num_5_index_1_share3, output_sum_secondmodule_equation_num_5_index_2_share3, output_sum_secondmodule_equation_num_5_index_3_share3, output_sum_secondmodule_equation_num_5_index_4_share3, output_sum_secondmodule_equation_num_5_index_5_share3, output_sum_secondmodule_equation_num_5_index_6_share3, output_sum_secondmodule_equation_num_5_index_7_share3, output_sum_secondmodule_equation_num_5_index_8_share3, output_sum_secondmodule_equation_num_5_index_9_share3, output_sum_secondmodule_equation_num_5_index_10_share3, output_sum_secondmodule_equation_num_5_index_11_share3, output_sum_secondmodule_equation_num_5_index_12_share3, output_sum_secondmodule_equation_num_5_index_13_share3, output_sum_secondmodule_equation_num_5_index_14_share3,
output_sum_secondmodule_equation_num_6_index_0_share3, output_sum_secondmodule_equation_num_6_index_1_share3, output_sum_secondmodule_equation_num_6_index_2_share3, output_sum_secondmodule_equation_num_6_index_3_share3, output_sum_secondmodule_equation_num_6_index_4_share3, output_sum_secondmodule_equation_num_6_index_5_share3, output_sum_secondmodule_equation_num_6_index_6_share3, output_sum_secondmodule_equation_num_6_index_7_share3, output_sum_secondmodule_equation_num_6_index_8_share3, output_sum_secondmodule_equation_num_6_index_9_share3, output_sum_secondmodule_equation_num_6_index_10_share3, output_sum_secondmodule_equation_num_6_index_11_share3, output_sum_secondmodule_equation_num_6_index_12_share3, output_sum_secondmodule_equation_num_6_index_13_share3, output_sum_secondmodule_equation_num_6_index_14_share3,
output_sum_secondmodule_equation_num_7_index_0_share3, output_sum_secondmodule_equation_num_7_index_1_share3, output_sum_secondmodule_equation_num_7_index_2_share3, output_sum_secondmodule_equation_num_7_index_3_share3, output_sum_secondmodule_equation_num_7_index_4_share3, output_sum_secondmodule_equation_num_7_index_5_share3, output_sum_secondmodule_equation_num_7_index_6_share3, output_sum_secondmodule_equation_num_7_index_7_share3, output_sum_secondmodule_equation_num_7_index_8_share3, output_sum_secondmodule_equation_num_7_index_9_share3, output_sum_secondmodule_equation_num_7_index_10_share3, output_sum_secondmodule_equation_num_7_index_11_share3, output_sum_secondmodule_equation_num_7_index_12_share3, output_sum_secondmodule_equation_num_7_index_13_share3, output_sum_secondmodule_equation_num_7_index_14_share3,
cross_module_equation_num0_domain_6, cross_module_equation_num1_domain_6, cross_module_equation_num2_domain_6, cross_module_equation_num3_domain_6,cross_module_equation_num4_domain_6,cross_module_equation_num5_domain_6,cross_module_equation_num6_domain_6,cross_module_equation_num7_domain_6
);



cross_module_multiplication inst_domain_7 (
output_x0_share3, output_x1_share3, output_x2_share3, output_x3_share3, output_x0x1_share3, output_x0x2_share3, output_x0x3_share3, output_x1x2_share3, output_x1x3_share3, output_x2x3_share3, output_x0x1x2_share3, output_x0x1x3_share3, output_x0x2x3_share3, output_x1x2x3_share3, output_x0x1x2x3_share3 , 
output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1,
cross_module_equation_num0_domain_7, cross_module_equation_num1_domain_7, cross_module_equation_num2_domain_7, cross_module_equation_num3_domain_7,cross_module_equation_num4_domain_7,cross_module_equation_num5_domain_7,cross_module_equation_num6_domain_7,cross_module_equation_num7_domain_7
);


cross_module_multiplication inst_domain_8 (
output_x0_share3, output_x1_share3, output_x2_share3, output_x3_share3, output_x0x1_share3, output_x0x2_share3, output_x0x3_share3, output_x1x2_share3, output_x1x3_share3, output_x2x3_share3, output_x0x1x2_share3, output_x0x1x3_share3, output_x0x2x3_share3, output_x1x2x3_share3, output_x0x1x2x3_share3 , 
output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2,
cross_module_equation_num0_domain_8, cross_module_equation_num1_domain_8, cross_module_equation_num2_domain_8, cross_module_equation_num3_domain_8,cross_module_equation_num4_domain_8,cross_module_equation_num5_domain_8,cross_module_equation_num6_domain_8,cross_module_equation_num7_domain_8
);


cross_module_multiplication inst_domain_9 (
output_x0_share3, output_x1_share3, output_x2_share3, output_x3_share3, output_x0x1_share3, output_x0x2_share3, output_x0x3_share3, output_x1x2_share3, output_x1x3_share3, output_x2x3_share3, output_x0x1x2_share3, output_x0x1x3_share3, output_x0x2x3_share3, output_x1x2x3_share3, output_x0x1x2x3_share3 , 
output_sum_secondmodule_equation_num_0_index_0_share3, output_sum_secondmodule_equation_num_0_index_1_share3, output_sum_secondmodule_equation_num_0_index_2_share3, output_sum_secondmodule_equation_num_0_index_3_share3, output_sum_secondmodule_equation_num_0_index_4_share3, output_sum_secondmodule_equation_num_0_index_5_share3, output_sum_secondmodule_equation_num_0_index_6_share3, output_sum_secondmodule_equation_num_0_index_7_share3, output_sum_secondmodule_equation_num_0_index_8_share3, output_sum_secondmodule_equation_num_0_index_9_share3, output_sum_secondmodule_equation_num_0_index_10_share3, output_sum_secondmodule_equation_num_0_index_11_share3, output_sum_secondmodule_equation_num_0_index_12_share3, output_sum_secondmodule_equation_num_0_index_13_share3, output_sum_secondmodule_equation_num_0_index_14_share3,
output_sum_secondmodule_equation_num_1_index_0_share3, output_sum_secondmodule_equation_num_1_index_1_share3, output_sum_secondmodule_equation_num_1_index_2_share3, output_sum_secondmodule_equation_num_1_index_3_share3, output_sum_secondmodule_equation_num_1_index_4_share3, output_sum_secondmodule_equation_num_1_index_5_share3, output_sum_secondmodule_equation_num_1_index_6_share3, output_sum_secondmodule_equation_num_1_index_7_share3, output_sum_secondmodule_equation_num_1_index_8_share3, output_sum_secondmodule_equation_num_1_index_9_share3, output_sum_secondmodule_equation_num_1_index_10_share3, output_sum_secondmodule_equation_num_1_index_11_share3, output_sum_secondmodule_equation_num_1_index_12_share3, output_sum_secondmodule_equation_num_1_index_13_share3, output_sum_secondmodule_equation_num_1_index_14_share3,
output_sum_secondmodule_equation_num_2_index_0_share3, output_sum_secondmodule_equation_num_2_index_1_share3, output_sum_secondmodule_equation_num_2_index_2_share3, output_sum_secondmodule_equation_num_2_index_3_share3, output_sum_secondmodule_equation_num_2_index_4_share3, output_sum_secondmodule_equation_num_2_index_5_share3, output_sum_secondmodule_equation_num_2_index_6_share3, output_sum_secondmodule_equation_num_2_index_7_share3, output_sum_secondmodule_equation_num_2_index_8_share3, output_sum_secondmodule_equation_num_2_index_9_share3, output_sum_secondmodule_equation_num_2_index_10_share3, output_sum_secondmodule_equation_num_2_index_11_share3, output_sum_secondmodule_equation_num_2_index_12_share3, output_sum_secondmodule_equation_num_2_index_13_share3, output_sum_secondmodule_equation_num_2_index_14_share3,
output_sum_secondmodule_equation_num_3_index_0_share3, output_sum_secondmodule_equation_num_3_index_1_share3, output_sum_secondmodule_equation_num_3_index_2_share3, output_sum_secondmodule_equation_num_3_index_3_share3, output_sum_secondmodule_equation_num_3_index_4_share3, output_sum_secondmodule_equation_num_3_index_5_share3, output_sum_secondmodule_equation_num_3_index_6_share3, output_sum_secondmodule_equation_num_3_index_7_share3, output_sum_secondmodule_equation_num_3_index_8_share3, output_sum_secondmodule_equation_num_3_index_9_share3, output_sum_secondmodule_equation_num_3_index_10_share3, output_sum_secondmodule_equation_num_3_index_11_share3, output_sum_secondmodule_equation_num_3_index_12_share3, output_sum_secondmodule_equation_num_3_index_13_share3, output_sum_secondmodule_equation_num_3_index_14_share3,
output_sum_secondmodule_equation_num_4_index_0_share3, output_sum_secondmodule_equation_num_4_index_1_share3, output_sum_secondmodule_equation_num_4_index_2_share3, output_sum_secondmodule_equation_num_4_index_3_share3, output_sum_secondmodule_equation_num_4_index_4_share3, output_sum_secondmodule_equation_num_4_index_5_share3, output_sum_secondmodule_equation_num_4_index_6_share3, output_sum_secondmodule_equation_num_4_index_7_share3, output_sum_secondmodule_equation_num_4_index_8_share3, output_sum_secondmodule_equation_num_4_index_9_share3, output_sum_secondmodule_equation_num_4_index_10_share3, output_sum_secondmodule_equation_num_4_index_11_share3, output_sum_secondmodule_equation_num_4_index_12_share3, output_sum_secondmodule_equation_num_4_index_13_share3, output_sum_secondmodule_equation_num_4_index_14_share3,
output_sum_secondmodule_equation_num_5_index_0_share3, output_sum_secondmodule_equation_num_5_index_1_share3, output_sum_secondmodule_equation_num_5_index_2_share3, output_sum_secondmodule_equation_num_5_index_3_share3, output_sum_secondmodule_equation_num_5_index_4_share3, output_sum_secondmodule_equation_num_5_index_5_share3, output_sum_secondmodule_equation_num_5_index_6_share3, output_sum_secondmodule_equation_num_5_index_7_share3, output_sum_secondmodule_equation_num_5_index_8_share3, output_sum_secondmodule_equation_num_5_index_9_share3, output_sum_secondmodule_equation_num_5_index_10_share3, output_sum_secondmodule_equation_num_5_index_11_share3, output_sum_secondmodule_equation_num_5_index_12_share3, output_sum_secondmodule_equation_num_5_index_13_share3, output_sum_secondmodule_equation_num_5_index_14_share3,
output_sum_secondmodule_equation_num_6_index_0_share3, output_sum_secondmodule_equation_num_6_index_1_share3, output_sum_secondmodule_equation_num_6_index_2_share3, output_sum_secondmodule_equation_num_6_index_3_share3, output_sum_secondmodule_equation_num_6_index_4_share3, output_sum_secondmodule_equation_num_6_index_5_share3, output_sum_secondmodule_equation_num_6_index_6_share3, output_sum_secondmodule_equation_num_6_index_7_share3, output_sum_secondmodule_equation_num_6_index_8_share3, output_sum_secondmodule_equation_num_6_index_9_share3, output_sum_secondmodule_equation_num_6_index_10_share3, output_sum_secondmodule_equation_num_6_index_11_share3, output_sum_secondmodule_equation_num_6_index_12_share3, output_sum_secondmodule_equation_num_6_index_13_share3, output_sum_secondmodule_equation_num_6_index_14_share3,
output_sum_secondmodule_equation_num_7_index_0_share3, output_sum_secondmodule_equation_num_7_index_1_share3, output_sum_secondmodule_equation_num_7_index_2_share3, output_sum_secondmodule_equation_num_7_index_3_share3, output_sum_secondmodule_equation_num_7_index_4_share3, output_sum_secondmodule_equation_num_7_index_5_share3, output_sum_secondmodule_equation_num_7_index_6_share3, output_sum_secondmodule_equation_num_7_index_7_share3, output_sum_secondmodule_equation_num_7_index_8_share3, output_sum_secondmodule_equation_num_7_index_9_share3, output_sum_secondmodule_equation_num_7_index_10_share3, output_sum_secondmodule_equation_num_7_index_11_share3, output_sum_secondmodule_equation_num_7_index_12_share3, output_sum_secondmodule_equation_num_7_index_13_share3, output_sum_secondmodule_equation_num_7_index_14_share3,
cross_module_equation_num0_domain_9, cross_module_equation_num1_domain_9, cross_module_equation_num2_domain_9, cross_module_equation_num3_domain_9,cross_module_equation_num4_domain_9,cross_module_equation_num5_domain_9,cross_module_equation_num6_domain_9,cross_module_equation_num7_domain_9
);


// Inner modules terms

first_and_second_inner domain_1_inst(   output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 ,   output_x4_share1, output_x5_share1, output_x6_share1, output_x7_share1, output_x4x5_share1, output_x4x6_share1, output_x4x7_share1, output_x5x6_share1, output_x5x7_share1, output_x6x7_share1, output_x4x5x6_share1, output_x4x5x7_share1, output_x4x6x7_share1, output_x5x6x7_share1, output_x4x5x6x7_share1 , inner_module_equation_num0_domain_1 , inner_module_equation_num1_domain_1 , inner_module_equation_num2_domain_1 , inner_module_equation_num3_domain_1 , inner_module_equation_num4_domain_1 , inner_module_equation_num5_domain_1 , inner_module_equation_num6_domain_1 , inner_module_equation_num7_domain_1 );

first_and_second_inner domain_5_inst(   output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 ,   output_x4_share2, output_x5_share2, output_x6_share2, output_x7_share2, output_x4x5_share2, output_x4x6_share2, output_x4x7_share2, output_x5x6_share2, output_x5x7_share2, output_x6x7_share2, output_x4x5x6_share2, output_x4x5x7_share2, output_x4x6x7_share2, output_x5x6x7_share2, output_x4x5x6x7_share2 , inner_module_equation_num0_domain_5 , inner_module_equation_num1_domain_5 , inner_module_equation_num2_domain_5 , inner_module_equation_num3_domain_5 , inner_module_equation_num4_domain_5 , inner_module_equation_num5_domain_5 , inner_module_equation_num6_domain_5 , inner_module_equation_num7_domain_5 );

first_and_second_inner domain_9_inst(   output_x0_share3, output_x1_share3, output_x2_share3, output_x3_share3, output_x0x1_share3, output_x0x2_share3, output_x0x3_share3, output_x1x2_share3, output_x1x3_share3, output_x2x3_share3, output_x0x1x2_share3, output_x0x1x3_share3, output_x0x2x3_share3, output_x1x2x3_share3, output_x0x1x2x3_share3 ,   output_x4_share3, output_x5_share3, output_x6_share3, output_x7_share3, output_x4x5_share3, output_x4x6_share3, output_x4x7_share3, output_x5x6_share3, output_x5x7_share3, output_x6x7_share3, output_x4x5x6_share3, output_x4x5x7_share3, output_x4x6x7_share3, output_x5x6x7_share3, output_x4x5x6x7_share3 , inner_module_equation_num0_domain_9 , inner_module_equation_num1_domain_9 , inner_module_equation_num2_domain_9 , inner_module_equation_num3_domain_9 , inner_module_equation_num4_domain_9 , inner_module_equation_num5_domain_9 , inner_module_equation_num6_domain_9 , inner_module_equation_num7_domain_9 );
 
wire inner_module_equation_num0_domain_2 ;
wire inner_module_equation_num1_domain_2 ;
wire inner_module_equation_num2_domain_2 ;
wire inner_module_equation_num3_domain_2 ;
wire inner_module_equation_num4_domain_2 ;
wire inner_module_equation_num5_domain_2 ;
wire inner_module_equation_num6_domain_2 ;
wire inner_module_equation_num7_domain_2 ;

assign inner_module_equation_num0_domain_2= 1'b0 ;
assign inner_module_equation_num1_domain_2= 1'b0 ;
assign inner_module_equation_num2_domain_2= 1'b0 ;
assign inner_module_equation_num3_domain_2= 1'b0 ;
assign inner_module_equation_num4_domain_2= 1'b0 ;
assign inner_module_equation_num5_domain_2= 1'b0 ;
assign inner_module_equation_num6_domain_2= 1'b0 ;
assign inner_module_equation_num7_domain_2= 1'b0 ;


wire inner_module_equation_num0_domain_3 ;
wire inner_module_equation_num1_domain_3 ;
wire inner_module_equation_num2_domain_3 ;
wire inner_module_equation_num3_domain_3 ;
wire inner_module_equation_num4_domain_3 ;
wire inner_module_equation_num5_domain_3 ;
wire inner_module_equation_num6_domain_3 ;
wire inner_module_equation_num7_domain_3 ;

assign inner_module_equation_num0_domain_3= 1'b0 ;
assign inner_module_equation_num1_domain_3= 1'b0 ;
assign inner_module_equation_num2_domain_3= 1'b0 ;
assign inner_module_equation_num3_domain_3= 1'b0 ;
assign inner_module_equation_num4_domain_3= 1'b0 ;
assign inner_module_equation_num5_domain_3= 1'b0 ;
assign inner_module_equation_num6_domain_3= 1'b0 ;
assign inner_module_equation_num7_domain_3= 1'b0 ;


wire inner_module_equation_num0_domain_4 ;
wire inner_module_equation_num1_domain_4 ;
wire inner_module_equation_num2_domain_4 ;
wire inner_module_equation_num3_domain_4 ;
wire inner_module_equation_num4_domain_4 ;
wire inner_module_equation_num5_domain_4 ;
wire inner_module_equation_num6_domain_4 ;
wire inner_module_equation_num7_domain_4 ;

assign inner_module_equation_num0_domain_4= 1'b0 ;
assign inner_module_equation_num1_domain_4= 1'b0 ;
assign inner_module_equation_num2_domain_4= 1'b0 ;
assign inner_module_equation_num3_domain_4= 1'b0 ;
assign inner_module_equation_num4_domain_4= 1'b0 ;
assign inner_module_equation_num5_domain_4= 1'b0 ;
assign inner_module_equation_num6_domain_4= 1'b0 ;
assign inner_module_equation_num7_domain_4= 1'b0 ;


wire inner_module_equation_num0_domain_6 ;
wire inner_module_equation_num1_domain_6 ;
wire inner_module_equation_num2_domain_6 ;
wire inner_module_equation_num3_domain_6 ;
wire inner_module_equation_num4_domain_6 ;
wire inner_module_equation_num5_domain_6 ;
wire inner_module_equation_num6_domain_6 ;
wire inner_module_equation_num7_domain_6 ;

assign inner_module_equation_num0_domain_6= 1'b0 ;
assign inner_module_equation_num1_domain_6= 1'b0 ;
assign inner_module_equation_num2_domain_6= 1'b0 ;
assign inner_module_equation_num3_domain_6= 1'b0 ;
assign inner_module_equation_num4_domain_6= 1'b0 ;
assign inner_module_equation_num5_domain_6= 1'b0 ;
assign inner_module_equation_num6_domain_6= 1'b0 ;
assign inner_module_equation_num7_domain_6= 1'b0 ;


wire inner_module_equation_num0_domain_7 ;
wire inner_module_equation_num1_domain_7 ;
wire inner_module_equation_num2_domain_7 ;
wire inner_module_equation_num3_domain_7 ;
wire inner_module_equation_num4_domain_7 ;
wire inner_module_equation_num5_domain_7 ;
wire inner_module_equation_num6_domain_7 ;
wire inner_module_equation_num7_domain_7 ;

assign inner_module_equation_num0_domain_7= 1'b0 ;
assign inner_module_equation_num1_domain_7= 1'b0 ;
assign inner_module_equation_num2_domain_7= 1'b0 ;
assign inner_module_equation_num3_domain_7= 1'b0 ;
assign inner_module_equation_num4_domain_7= 1'b0 ;
assign inner_module_equation_num5_domain_7= 1'b0 ;
assign inner_module_equation_num6_domain_7= 1'b0 ;
assign inner_module_equation_num7_domain_7= 1'b0 ;


wire inner_module_equation_num0_domain_8 ;
wire inner_module_equation_num1_domain_8 ;
wire inner_module_equation_num2_domain_8 ;
wire inner_module_equation_num3_domain_8 ;
wire inner_module_equation_num4_domain_8 ;
wire inner_module_equation_num5_domain_8 ;
wire inner_module_equation_num6_domain_8 ;
wire inner_module_equation_num7_domain_8 ;

assign inner_module_equation_num0_domain_8= 1'b0 ;
assign inner_module_equation_num1_domain_8= 1'b0 ;
assign inner_module_equation_num2_domain_8= 1'b0 ;
assign inner_module_equation_num3_domain_8= 1'b0 ;
assign inner_module_equation_num4_domain_8= 1'b0 ;
assign inner_module_equation_num5_domain_8= 1'b0 ;
assign inner_module_equation_num6_domain_8= 1'b0 ;
assign inner_module_equation_num7_domain_8= 1'b0 ;


// Merge inner and cross domains

xor_module xor_num0_dom1(cross_module_equation_num0_domain_1,inner_module_equation_num0_domain_1,inner_plus_cross_module_equation_num0_domain_1);
xor_module xor_num0_dom2(cross_module_equation_num0_domain_2,inner_module_equation_num0_domain_2,inner_plus_cross_module_equation_num0_domain_2);
xor_module xor_num0_dom3(cross_module_equation_num0_domain_3,inner_module_equation_num0_domain_3,inner_plus_cross_module_equation_num0_domain_3);
xor_module xor_num0_dom4(cross_module_equation_num0_domain_4,inner_module_equation_num0_domain_4,inner_plus_cross_module_equation_num0_domain_4);
xor_module xor_num0_dom5(cross_module_equation_num0_domain_5,inner_module_equation_num0_domain_5,inner_plus_cross_module_equation_num0_domain_5);
xor_module xor_num0_dom6(cross_module_equation_num0_domain_6,inner_module_equation_num0_domain_6,inner_plus_cross_module_equation_num0_domain_6);
xor_module xor_num0_dom7(cross_module_equation_num0_domain_7,inner_module_equation_num0_domain_7,inner_plus_cross_module_equation_num0_domain_7);
xor_module xor_num0_dom8(cross_module_equation_num0_domain_8,inner_module_equation_num0_domain_8,inner_plus_cross_module_equation_num0_domain_8);
xor_module xor_num0_dom9(cross_module_equation_num0_domain_9,inner_module_equation_num0_domain_9,inner_plus_cross_module_equation_num0_domain_9);



xor_module xor_num1_dom1(cross_module_equation_num1_domain_1,inner_module_equation_num1_domain_1,inner_plus_cross_module_equation_num1_domain_1);
xor_module xor_num1_dom2(cross_module_equation_num1_domain_2,inner_module_equation_num1_domain_2,inner_plus_cross_module_equation_num1_domain_2);
xor_module xor_num1_dom3(cross_module_equation_num1_domain_3,inner_module_equation_num1_domain_3,inner_plus_cross_module_equation_num1_domain_3);
xor_module xor_num1_dom4(cross_module_equation_num1_domain_4,inner_module_equation_num1_domain_4,inner_plus_cross_module_equation_num1_domain_4);
xor_module xor_num1_dom5(cross_module_equation_num1_domain_5,inner_module_equation_num1_domain_5,inner_plus_cross_module_equation_num1_domain_5);
xor_module xor_num1_dom6(cross_module_equation_num1_domain_6,inner_module_equation_num1_domain_6,inner_plus_cross_module_equation_num1_domain_6);
xor_module xor_num1_dom7(cross_module_equation_num1_domain_7,inner_module_equation_num1_domain_7,inner_plus_cross_module_equation_num1_domain_7);
xor_module xor_num1_dom8(cross_module_equation_num1_domain_8,inner_module_equation_num1_domain_8,inner_plus_cross_module_equation_num1_domain_8);
xor_module xor_num1_dom9(cross_module_equation_num1_domain_9,inner_module_equation_num1_domain_9,inner_plus_cross_module_equation_num1_domain_9);



xor_module xor_num2_dom1(cross_module_equation_num2_domain_1,inner_module_equation_num2_domain_1,inner_plus_cross_module_equation_num2_domain_1);
xor_module xor_num2_dom2(cross_module_equation_num2_domain_2,inner_module_equation_num2_domain_2,inner_plus_cross_module_equation_num2_domain_2);
xor_module xor_num2_dom3(cross_module_equation_num2_domain_3,inner_module_equation_num2_domain_3,inner_plus_cross_module_equation_num2_domain_3);
xor_module xor_num2_dom4(cross_module_equation_num2_domain_4,inner_module_equation_num2_domain_4,inner_plus_cross_module_equation_num2_domain_4);
xor_module xor_num2_dom5(cross_module_equation_num2_domain_5,inner_module_equation_num2_domain_5,inner_plus_cross_module_equation_num2_domain_5);
xor_module xor_num2_dom6(cross_module_equation_num2_domain_6,inner_module_equation_num2_domain_6,inner_plus_cross_module_equation_num2_domain_6);
xor_module xor_num2_dom7(cross_module_equation_num2_domain_7,inner_module_equation_num2_domain_7,inner_plus_cross_module_equation_num2_domain_7);
xor_module xor_num2_dom8(cross_module_equation_num2_domain_8,inner_module_equation_num2_domain_8,inner_plus_cross_module_equation_num2_domain_8);
xor_module xor_num2_dom9(cross_module_equation_num2_domain_9,inner_module_equation_num2_domain_9,inner_plus_cross_module_equation_num2_domain_9);



xor_module xor_num3_dom1(cross_module_equation_num3_domain_1,inner_module_equation_num3_domain_1,inner_plus_cross_module_equation_num3_domain_1);
xor_module xor_num3_dom2(cross_module_equation_num3_domain_2,inner_module_equation_num3_domain_2,inner_plus_cross_module_equation_num3_domain_2);
xor_module xor_num3_dom3(cross_module_equation_num3_domain_3,inner_module_equation_num3_domain_3,inner_plus_cross_module_equation_num3_domain_3);
xor_module xor_num3_dom4(cross_module_equation_num3_domain_4,inner_module_equation_num3_domain_4,inner_plus_cross_module_equation_num3_domain_4);
xor_module xor_num3_dom5(cross_module_equation_num3_domain_5,inner_module_equation_num3_domain_5,inner_plus_cross_module_equation_num3_domain_5);
xor_module xor_num3_dom6(cross_module_equation_num3_domain_6,inner_module_equation_num3_domain_6,inner_plus_cross_module_equation_num3_domain_6);
xor_module xor_num3_dom7(cross_module_equation_num3_domain_7,inner_module_equation_num3_domain_7,inner_plus_cross_module_equation_num3_domain_7);
xor_module xor_num3_dom8(cross_module_equation_num3_domain_8,inner_module_equation_num3_domain_8,inner_plus_cross_module_equation_num3_domain_8);
xor_module xor_num3_dom9(cross_module_equation_num3_domain_9,inner_module_equation_num3_domain_9,inner_plus_cross_module_equation_num3_domain_9);



xor_module xor_num4_dom1(cross_module_equation_num4_domain_1,inner_module_equation_num4_domain_1,inner_plus_cross_module_equation_num4_domain_1);
xor_module xor_num4_dom2(cross_module_equation_num4_domain_2,inner_module_equation_num4_domain_2,inner_plus_cross_module_equation_num4_domain_2);
xor_module xor_num4_dom3(cross_module_equation_num4_domain_3,inner_module_equation_num4_domain_3,inner_plus_cross_module_equation_num4_domain_3);
xor_module xor_num4_dom4(cross_module_equation_num4_domain_4,inner_module_equation_num4_domain_4,inner_plus_cross_module_equation_num4_domain_4);
xor_module xor_num4_dom5(cross_module_equation_num4_domain_5,inner_module_equation_num4_domain_5,inner_plus_cross_module_equation_num4_domain_5);
xor_module xor_num4_dom6(cross_module_equation_num4_domain_6,inner_module_equation_num4_domain_6,inner_plus_cross_module_equation_num4_domain_6);
xor_module xor_num4_dom7(cross_module_equation_num4_domain_7,inner_module_equation_num4_domain_7,inner_plus_cross_module_equation_num4_domain_7);
xor_module xor_num4_dom8(cross_module_equation_num4_domain_8,inner_module_equation_num4_domain_8,inner_plus_cross_module_equation_num4_domain_8);
xor_module xor_num4_dom9(cross_module_equation_num4_domain_9,inner_module_equation_num4_domain_9,inner_plus_cross_module_equation_num4_domain_9);


xor_module xor_num5_dom1(cross_module_equation_num5_domain_1,inner_module_equation_num5_domain_1,inner_plus_cross_module_equation_num5_domain_1);
xor_module xor_num5_dom2(cross_module_equation_num5_domain_2,inner_module_equation_num5_domain_2,inner_plus_cross_module_equation_num5_domain_2);
xor_module xor_num5_dom3(cross_module_equation_num5_domain_3,inner_module_equation_num5_domain_3,inner_plus_cross_module_equation_num5_domain_3);
xor_module xor_num5_dom4(cross_module_equation_num5_domain_4,inner_module_equation_num5_domain_4,inner_plus_cross_module_equation_num5_domain_4);
xor_module xor_num5_dom5(cross_module_equation_num5_domain_5,inner_module_equation_num5_domain_5,inner_plus_cross_module_equation_num5_domain_5);
xor_module xor_num5_dom6(cross_module_equation_num5_domain_6,inner_module_equation_num5_domain_6,inner_plus_cross_module_equation_num5_domain_6);
xor_module xor_num5_dom7(cross_module_equation_num5_domain_7,inner_module_equation_num5_domain_7,inner_plus_cross_module_equation_num5_domain_7);
xor_module xor_num5_dom8(cross_module_equation_num5_domain_8,inner_module_equation_num5_domain_8,inner_plus_cross_module_equation_num5_domain_8);
xor_module xor_num5_dom9(cross_module_equation_num5_domain_9,inner_module_equation_num5_domain_9,inner_plus_cross_module_equation_num5_domain_9);


xor_module xor_num6_dom1(cross_module_equation_num6_domain_1,inner_module_equation_num6_domain_1,inner_plus_cross_module_equation_num6_domain_1);
xor_module xor_num6_dom2(cross_module_equation_num6_domain_2,inner_module_equation_num6_domain_2,inner_plus_cross_module_equation_num6_domain_2);
xor_module xor_num6_dom3(cross_module_equation_num6_domain_3,inner_module_equation_num6_domain_3,inner_plus_cross_module_equation_num6_domain_3);
xor_module xor_num6_dom4(cross_module_equation_num6_domain_4,inner_module_equation_num6_domain_4,inner_plus_cross_module_equation_num6_domain_4);
xor_module xor_num6_dom5(cross_module_equation_num6_domain_5,inner_module_equation_num6_domain_5,inner_plus_cross_module_equation_num6_domain_5);
xor_module xor_num6_dom6(cross_module_equation_num6_domain_6,inner_module_equation_num6_domain_6,inner_plus_cross_module_equation_num6_domain_6);
xor_module xor_num6_dom7(cross_module_equation_num6_domain_7,inner_module_equation_num6_domain_7,inner_plus_cross_module_equation_num6_domain_7);
xor_module xor_num6_dom8(cross_module_equation_num6_domain_8,inner_module_equation_num6_domain_8,inner_plus_cross_module_equation_num6_domain_8);
xor_module xor_num6_dom9(cross_module_equation_num6_domain_9,inner_module_equation_num6_domain_9,inner_plus_cross_module_equation_num6_domain_9);


xor_module xor_num7_dom1(cross_module_equation_num7_domain_1,inner_module_equation_num7_domain_1,inner_plus_cross_module_equation_num7_domain_1);
xor_module xor_num7_dom2(cross_module_equation_num7_domain_2,inner_module_equation_num7_domain_2,inner_plus_cross_module_equation_num7_domain_2);
xor_module xor_num7_dom3(cross_module_equation_num7_domain_3,inner_module_equation_num7_domain_3,inner_plus_cross_module_equation_num7_domain_3);
xor_module xor_num7_dom4(cross_module_equation_num7_domain_4,inner_module_equation_num7_domain_4,inner_plus_cross_module_equation_num7_domain_4);
xor_module xor_num7_dom5(cross_module_equation_num7_domain_5,inner_module_equation_num7_domain_5,inner_plus_cross_module_equation_num7_domain_5);
xor_module xor_num7_dom6(cross_module_equation_num7_domain_6,inner_module_equation_num7_domain_6,inner_plus_cross_module_equation_num7_domain_6);
xor_module xor_num7_dom7(cross_module_equation_num7_domain_7,inner_module_equation_num7_domain_7,inner_plus_cross_module_equation_num7_domain_7);
xor_module xor_num7_dom8(cross_module_equation_num7_domain_8,inner_module_equation_num7_domain_8,inner_plus_cross_module_equation_num7_domain_8);
xor_module xor_num7_dom9(cross_module_equation_num7_domain_9,inner_module_equation_num7_domain_9,inner_plus_cross_module_equation_num7_domain_9);


// Refresh and store in registers

wire [3:1] rand_bit_num0, rand_bit_num1, rand_bit_num2, rand_bit_num3, rand_bit_num4, rand_bit_num5, rand_bit_num6, rand_bit_num7;
assign rand_bit_num0 = rand_bit_second[3:1];
assign rand_bit_num1 = rand_bit_second[6:4];
assign rand_bit_num2 = rand_bit_second[9:7];
assign rand_bit_num3 = rand_bit_second[12:10];
assign rand_bit_num4 = rand_bit_second[15:13];
assign rand_bit_num5 = rand_bit_second[18:16];
assign rand_bit_num6 = rand_bit_second[21:19];
assign rand_bit_num7 = rand_bit_second[24:22];

reg sbox_out_num0_domain_1_reg,sbox_out_num0_domain_2_reg,sbox_out_num0_domain_3_reg, sbox_out_num0_domain_4_reg, sbox_out_num0_domain_5_reg, sbox_out_num0_domain_6_reg, sbox_out_num0_domain_7_reg, sbox_out_num0_domain_8_reg, sbox_out_num0_domain_9_reg;

always@(posedge clk)
begin
        sbox_out_num0_domain_1_reg <= inner_plus_cross_module_equation_num0_domain_1 ^ 1'b1;
        sbox_out_num0_domain_2_reg <= inner_plus_cross_module_equation_num0_domain_2 ^ rand_bit_num0[1];
        sbox_out_num0_domain_3_reg <= inner_plus_cross_module_equation_num0_domain_3 ^ rand_bit_num0[2];
        sbox_out_num0_domain_4_reg <= inner_plus_cross_module_equation_num0_domain_4 ^ rand_bit_num0[1];
        sbox_out_num0_domain_5_reg <= inner_plus_cross_module_equation_num0_domain_5 ;
        sbox_out_num0_domain_6_reg <= inner_plus_cross_module_equation_num0_domain_6 ^ rand_bit_num0[3];
        sbox_out_num0_domain_7_reg <= inner_plus_cross_module_equation_num0_domain_7 ^ rand_bit_num0[2];
        sbox_out_num0_domain_8_reg <= inner_plus_cross_module_equation_num0_domain_8 ^ rand_bit_num0[3];
        sbox_out_num0_domain_9_reg <= inner_plus_cross_module_equation_num0_domain_9 ;
end

wire sbox_out_num0_share1, sbox_out_num0_share2 , sbox_out_num0_share3 ;
assign sbox_out_num0_share1 = sbox_out_num0_domain_1_reg ^ sbox_out_num0_domain_2_reg ^ sbox_out_num0_domain_3_reg ;
assign sbox_out_num0_share2 = sbox_out_num0_domain_4_reg ^ sbox_out_num0_domain_5_reg ^ sbox_out_num0_domain_6_reg ;
assign sbox_out_num0_share3 = sbox_out_num0_domain_7_reg ^ sbox_out_num0_domain_8_reg ^ sbox_out_num0_domain_9_reg ;




reg sbox_out_num1_domain_1_reg,sbox_out_num1_domain_2_reg,sbox_out_num1_domain_3_reg, sbox_out_num1_domain_4_reg, sbox_out_num1_domain_5_reg, sbox_out_num1_domain_6_reg, sbox_out_num1_domain_7_reg, sbox_out_num1_domain_8_reg, sbox_out_num1_domain_9_reg;

always@(posedge clk)
begin
        sbox_out_num1_domain_1_reg <= inner_plus_cross_module_equation_num1_domain_1 ^ 1'b1;
        sbox_out_num1_domain_2_reg <= inner_plus_cross_module_equation_num1_domain_2 ^ rand_bit_num1[1];
        sbox_out_num1_domain_3_reg <= inner_plus_cross_module_equation_num1_domain_3 ^ rand_bit_num1[2];
        sbox_out_num1_domain_4_reg <= inner_plus_cross_module_equation_num1_domain_4 ^ rand_bit_num1[1];
        sbox_out_num1_domain_5_reg <= inner_plus_cross_module_equation_num1_domain_5 ;
        sbox_out_num1_domain_6_reg <= inner_plus_cross_module_equation_num1_domain_6 ^ rand_bit_num1[3];
        sbox_out_num1_domain_7_reg <= inner_plus_cross_module_equation_num1_domain_7 ^ rand_bit_num1[2];
        sbox_out_num1_domain_8_reg <= inner_plus_cross_module_equation_num1_domain_8 ^ rand_bit_num1[3];
        sbox_out_num1_domain_9_reg <= inner_plus_cross_module_equation_num1_domain_9 ;
end

wire sbox_out_num1_share1, sbox_out_num1_share2 , sbox_out_num1_share3 ;
assign sbox_out_num1_share1 = sbox_out_num1_domain_1_reg ^ sbox_out_num1_domain_2_reg ^ sbox_out_num1_domain_3_reg ;
assign sbox_out_num1_share2 = sbox_out_num1_domain_4_reg ^ sbox_out_num1_domain_5_reg ^ sbox_out_num1_domain_6_reg ;
assign sbox_out_num1_share3 = sbox_out_num1_domain_7_reg ^ sbox_out_num1_domain_8_reg ^ sbox_out_num1_domain_9_reg ;





reg sbox_out_num2_domain_1_reg,sbox_out_num2_domain_2_reg,sbox_out_num2_domain_3_reg, sbox_out_num2_domain_4_reg, sbox_out_num2_domain_5_reg, sbox_out_num2_domain_6_reg, sbox_out_num2_domain_7_reg, sbox_out_num2_domain_8_reg, sbox_out_num2_domain_9_reg;

always@(posedge clk)
begin
        sbox_out_num2_domain_1_reg <= inner_plus_cross_module_equation_num2_domain_1 ;
        sbox_out_num2_domain_2_reg <= inner_plus_cross_module_equation_num2_domain_2 ^ rand_bit_num2[1];
        sbox_out_num2_domain_3_reg <= inner_plus_cross_module_equation_num2_domain_3 ^ rand_bit_num2[2];
        sbox_out_num2_domain_4_reg <= inner_plus_cross_module_equation_num2_domain_4 ^ rand_bit_num2[1];
        sbox_out_num2_domain_5_reg <= inner_plus_cross_module_equation_num2_domain_5 ;
        sbox_out_num2_domain_6_reg <= inner_plus_cross_module_equation_num2_domain_6 ^ rand_bit_num2[3];
        sbox_out_num2_domain_7_reg <= inner_plus_cross_module_equation_num2_domain_7 ^ rand_bit_num2[2];
        sbox_out_num2_domain_8_reg <= inner_plus_cross_module_equation_num2_domain_8 ^ rand_bit_num2[3];
        sbox_out_num2_domain_9_reg <= inner_plus_cross_module_equation_num2_domain_9 ;
end

wire sbox_out_num2_share1, sbox_out_num2_share2 , sbox_out_num2_share3 ;
assign sbox_out_num2_share1 = sbox_out_num2_domain_1_reg ^ sbox_out_num2_domain_2_reg ^ sbox_out_num2_domain_3_reg ;
assign sbox_out_num2_share2 = sbox_out_num2_domain_4_reg ^ sbox_out_num2_domain_5_reg ^ sbox_out_num2_domain_6_reg ;
assign sbox_out_num2_share3 = sbox_out_num2_domain_7_reg ^ sbox_out_num2_domain_8_reg ^ sbox_out_num2_domain_9_reg ;




reg sbox_out_num3_domain_1_reg,sbox_out_num3_domain_2_reg,sbox_out_num3_domain_3_reg, sbox_out_num3_domain_4_reg, sbox_out_num3_domain_5_reg, sbox_out_num3_domain_6_reg, sbox_out_num3_domain_7_reg, sbox_out_num3_domain_8_reg, sbox_out_num3_domain_9_reg;

always@(posedge clk)
begin
        sbox_out_num3_domain_1_reg <= inner_plus_cross_module_equation_num3_domain_1 ;
        sbox_out_num3_domain_2_reg <= inner_plus_cross_module_equation_num3_domain_2 ^ rand_bit_num3[1];
        sbox_out_num3_domain_3_reg <= inner_plus_cross_module_equation_num3_domain_3 ^ rand_bit_num3[2];
        sbox_out_num3_domain_4_reg <= inner_plus_cross_module_equation_num3_domain_4 ^ rand_bit_num3[1];
        sbox_out_num3_domain_5_reg <= inner_plus_cross_module_equation_num3_domain_5 ;
        sbox_out_num3_domain_6_reg <= inner_plus_cross_module_equation_num3_domain_6 ^ rand_bit_num3[3];
        sbox_out_num3_domain_7_reg <= inner_plus_cross_module_equation_num3_domain_7 ^ rand_bit_num3[2];
        sbox_out_num3_domain_8_reg <= inner_plus_cross_module_equation_num3_domain_8 ^ rand_bit_num3[3];
        sbox_out_num3_domain_9_reg <= inner_plus_cross_module_equation_num3_domain_9 ;
end

wire sbox_out_num3_share1, sbox_out_num3_share2 , sbox_out_num3_share3 ;
assign sbox_out_num3_share1 = sbox_out_num3_domain_1_reg ^ sbox_out_num3_domain_2_reg ^ sbox_out_num3_domain_3_reg ;
assign sbox_out_num3_share2 = sbox_out_num3_domain_4_reg ^ sbox_out_num3_domain_5_reg ^ sbox_out_num3_domain_6_reg ;
assign sbox_out_num3_share3 = sbox_out_num3_domain_7_reg ^ sbox_out_num3_domain_8_reg ^ sbox_out_num3_domain_9_reg ;


reg sbox_out_num4_domain_1_reg,sbox_out_num4_domain_2_reg,sbox_out_num4_domain_3_reg, sbox_out_num4_domain_4_reg, sbox_out_num4_domain_5_reg, sbox_out_num4_domain_6_reg, sbox_out_num4_domain_7_reg, sbox_out_num4_domain_8_reg, sbox_out_num4_domain_9_reg;

always@(posedge clk)
begin
        sbox_out_num4_domain_1_reg <= inner_plus_cross_module_equation_num4_domain_1 ;
        sbox_out_num4_domain_2_reg <= inner_plus_cross_module_equation_num4_domain_2 ^ rand_bit_num4[1];
        sbox_out_num4_domain_3_reg <= inner_plus_cross_module_equation_num4_domain_3 ^ rand_bit_num4[2];
        sbox_out_num4_domain_4_reg <= inner_plus_cross_module_equation_num4_domain_4 ^ rand_bit_num4[1];
        sbox_out_num4_domain_5_reg <= inner_plus_cross_module_equation_num4_domain_5 ;
        sbox_out_num4_domain_6_reg <= inner_plus_cross_module_equation_num4_domain_6 ^ rand_bit_num4[3];
        sbox_out_num4_domain_7_reg <= inner_plus_cross_module_equation_num4_domain_7 ^ rand_bit_num4[2];
        sbox_out_num4_domain_8_reg <= inner_plus_cross_module_equation_num4_domain_8 ^ rand_bit_num4[3];
        sbox_out_num4_domain_9_reg <= inner_plus_cross_module_equation_num4_domain_9 ;
end

wire sbox_out_num4_share1, sbox_out_num4_share2 , sbox_out_num4_share3 ;
assign sbox_out_num4_share1 = sbox_out_num4_domain_1_reg ^ sbox_out_num4_domain_2_reg ^ sbox_out_num4_domain_3_reg ;
assign sbox_out_num4_share2 = sbox_out_num4_domain_4_reg ^ sbox_out_num4_domain_5_reg ^ sbox_out_num4_domain_6_reg ;
assign sbox_out_num4_share3 = sbox_out_num4_domain_7_reg ^ sbox_out_num4_domain_8_reg ^ sbox_out_num4_domain_9_reg ;




reg sbox_out_num5_domain_1_reg,sbox_out_num5_domain_2_reg,sbox_out_num5_domain_3_reg, sbox_out_num5_domain_4_reg, sbox_out_num5_domain_5_reg, sbox_out_num5_domain_6_reg, sbox_out_num5_domain_7_reg, sbox_out_num5_domain_8_reg, sbox_out_num5_domain_9_reg;

always@(posedge clk)
begin
        sbox_out_num5_domain_1_reg <= inner_plus_cross_module_equation_num5_domain_1 ^ 1'b1;
        sbox_out_num5_domain_2_reg <= inner_plus_cross_module_equation_num5_domain_2 ^ rand_bit_num5[1];
        sbox_out_num5_domain_3_reg <= inner_plus_cross_module_equation_num5_domain_3 ^ rand_bit_num5[2];
        sbox_out_num5_domain_4_reg <= inner_plus_cross_module_equation_num5_domain_4 ^ rand_bit_num5[1];
        sbox_out_num5_domain_5_reg <= inner_plus_cross_module_equation_num5_domain_5 ;
        sbox_out_num5_domain_6_reg <= inner_plus_cross_module_equation_num5_domain_6 ^ rand_bit_num5[3];
        sbox_out_num5_domain_7_reg <= inner_plus_cross_module_equation_num5_domain_7 ^ rand_bit_num5[2];
        sbox_out_num5_domain_8_reg <= inner_plus_cross_module_equation_num5_domain_8 ^ rand_bit_num5[3];
        sbox_out_num5_domain_9_reg <= inner_plus_cross_module_equation_num5_domain_9 ;
end

wire sbox_out_num5_share1, sbox_out_num5_share2 , sbox_out_num5_share3 ;
assign sbox_out_num5_share1 = sbox_out_num5_domain_1_reg ^ sbox_out_num5_domain_2_reg ^ sbox_out_num5_domain_3_reg ;
assign sbox_out_num5_share2 = sbox_out_num5_domain_4_reg ^ sbox_out_num5_domain_5_reg ^ sbox_out_num5_domain_6_reg ;
assign sbox_out_num5_share3 = sbox_out_num5_domain_7_reg ^ sbox_out_num5_domain_8_reg ^ sbox_out_num5_domain_9_reg ;



reg sbox_out_num6_domain_1_reg,sbox_out_num6_domain_2_reg,sbox_out_num6_domain_3_reg, sbox_out_num6_domain_4_reg, sbox_out_num6_domain_5_reg, sbox_out_num6_domain_6_reg, sbox_out_num6_domain_7_reg, sbox_out_num6_domain_8_reg, sbox_out_num6_domain_9_reg;

always@(posedge clk)
begin
        sbox_out_num6_domain_1_reg <= inner_plus_cross_module_equation_num6_domain_1 ^ 1'b1;
        sbox_out_num6_domain_2_reg <= inner_plus_cross_module_equation_num6_domain_2 ^ rand_bit_num6[1];
        sbox_out_num6_domain_3_reg <= inner_plus_cross_module_equation_num6_domain_3 ^ rand_bit_num6[2];
        sbox_out_num6_domain_4_reg <= inner_plus_cross_module_equation_num6_domain_4 ^ rand_bit_num6[1];
        sbox_out_num6_domain_5_reg <= inner_plus_cross_module_equation_num6_domain_5 ;
        sbox_out_num6_domain_6_reg <= inner_plus_cross_module_equation_num6_domain_6 ^ rand_bit_num6[3];
        sbox_out_num6_domain_7_reg <= inner_plus_cross_module_equation_num6_domain_7 ^ rand_bit_num6[2];
        sbox_out_num6_domain_8_reg <= inner_plus_cross_module_equation_num6_domain_8 ^ rand_bit_num6[3];
        sbox_out_num6_domain_9_reg <= inner_plus_cross_module_equation_num6_domain_9 ;
end

wire sbox_out_num6_share1, sbox_out_num6_share2 , sbox_out_num6_share3 ;
assign sbox_out_num6_share1 = sbox_out_num6_domain_1_reg ^ sbox_out_num6_domain_2_reg ^ sbox_out_num6_domain_3_reg ;
assign sbox_out_num6_share2 = sbox_out_num6_domain_4_reg ^ sbox_out_num6_domain_5_reg ^ sbox_out_num6_domain_6_reg ;
assign sbox_out_num6_share3 = sbox_out_num6_domain_7_reg ^ sbox_out_num6_domain_8_reg ^ sbox_out_num6_domain_9_reg ;



reg sbox_out_num7_domain_1_reg,sbox_out_num7_domain_2_reg,sbox_out_num7_domain_3_reg, sbox_out_num7_domain_4_reg, sbox_out_num7_domain_5_reg, sbox_out_num7_domain_6_reg, sbox_out_num7_domain_7_reg, sbox_out_num7_domain_8_reg, sbox_out_num7_domain_9_reg;

always@(posedge clk)
begin
        sbox_out_num7_domain_1_reg <= inner_plus_cross_module_equation_num7_domain_1 ;
        sbox_out_num7_domain_2_reg <= inner_plus_cross_module_equation_num7_domain_2 ^ rand_bit_num7[1];
        sbox_out_num7_domain_3_reg <= inner_plus_cross_module_equation_num7_domain_3 ^ rand_bit_num7[2];
        sbox_out_num7_domain_4_reg <= inner_plus_cross_module_equation_num7_domain_4 ^ rand_bit_num7[1];
        sbox_out_num7_domain_5_reg <= inner_plus_cross_module_equation_num7_domain_5 ;
        sbox_out_num7_domain_6_reg <= inner_plus_cross_module_equation_num7_domain_6 ^ rand_bit_num7[3];
        sbox_out_num7_domain_7_reg <= inner_plus_cross_module_equation_num7_domain_7 ^ rand_bit_num7[2];
        sbox_out_num7_domain_8_reg <= inner_plus_cross_module_equation_num7_domain_8 ^ rand_bit_num7[3];
        sbox_out_num7_domain_9_reg <= inner_plus_cross_module_equation_num7_domain_9 ;
end

wire sbox_out_num7_share1, sbox_out_num7_share2 , sbox_out_num7_share3 ;
assign sbox_out_num7_share1 = sbox_out_num7_domain_1_reg ^ sbox_out_num7_domain_2_reg ^ sbox_out_num7_domain_3_reg ;
assign sbox_out_num7_share2 = sbox_out_num7_domain_4_reg ^ sbox_out_num7_domain_5_reg ^ sbox_out_num7_domain_6_reg ;
assign sbox_out_num7_share3 = sbox_out_num7_domain_7_reg ^ sbox_out_num7_domain_8_reg ^ sbox_out_num7_domain_9_reg ;



// Assign outputs


assign output_sbox_share1 = {sbox_out_num7_share1,sbox_out_num6_share1,sbox_out_num5_share1,sbox_out_num4_share1,sbox_out_num3_share1,sbox_out_num2_share1,sbox_out_num1_share1,sbox_out_num0_share1};
assign output_sbox_share2 = {sbox_out_num7_share2,sbox_out_num6_share2,sbox_out_num5_share2,sbox_out_num4_share2,sbox_out_num3_share2,sbox_out_num2_share2,sbox_out_num1_share2,sbox_out_num0_share2};
assign output_sbox_share3 = {sbox_out_num7_share3,sbox_out_num6_share3,sbox_out_num5_share3,sbox_out_num4_share3,sbox_out_num3_share3,sbox_out_num2_share3,sbox_out_num1_share3,sbox_out_num0_share3};

endmodule