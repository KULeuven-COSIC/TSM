`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 22:00:00 02/22/2025
// Design Name: XOR Operation for One Share
// Module Name: xor_AES_twofiftyfour
// Project Name: AES Masked S-Box
// Target Device: FPGA
// Tool Versions: Vivado 2020.2
// Description: Computes bitwise XOR of 254 input signals for exactly one share.
// Dependencies: None
//
// Revision:
// Revision 0.01 - Initial version
//
//////////////////////////////////////////////////////////////////////////////////


module xor_AES_twofiftyfour(
in1_1 , in1_2 , in1_3 , in1_4 , in1_5 , in1_6 , in1_7 , in1_8 , in1_9 , in1_10 , in1_11 , in1_12 , in1_13 , in1_14 , in1_15 , in1_16 , in1_17 , in1_18 , in1_19 , in1_20 , in1_21 , in1_22 , in1_23 , in1_24 , in1_25 , in1_26 , in1_27 , in1_28 , in1_29 , in1_30 , in1_31 , in1_32 , in1_33 , in1_34 , in1_35 , in1_36 , in1_37 , in1_38 , in1_39 , in1_40 , in1_41 , in1_42 , in1_43 , in1_44 , in1_45 , in1_46 , in1_47 , in1_48 , in1_49 , in1_50 , in1_51 , in1_52 , in1_53 , in1_54 , in1_55 , in1_56 , in1_57 , in1_58 , in1_59 , in1_60 , in1_61 , in1_62 , in1_63 , in1_64 , in1_65 , in1_66 , in1_67 , in1_68 , in1_69 , in1_70 , in1_71 , in1_72 , in1_73 , in1_74 , in1_75 , in1_76 , in1_77 , in1_78 , in1_79 , in1_80 , in1_81 , in1_82 , in1_83 , in1_84 , in1_85 , in1_86 , in1_87 , in1_88 , in1_89 , in1_90 , in1_91 , in1_92 , in1_93 , in1_94 , in1_95 , in1_96 , in1_97 , in1_98 , in1_99 , in1_100 , in1_101 , in1_102 , in1_103 , in1_104 , in1_105 , in1_106 , in1_107 , in1_108 , in1_109 , in1_110 , in1_111 , in1_112 , in1_113 , in1_114 , in1_115 , in1_116 , in1_117 , in1_118 , in1_119 , in1_120 , in1_121 , in1_122 , in1_123 , in1_124 , in1_125 , in1_126 , in1_127 , in1_128 , in1_129 , in1_130 , in1_131 , in1_132 , in1_133 , in1_134 , in1_135 , in1_136 , in1_137 , in1_138 , in1_139 , in1_140 , in1_141 , in1_142 , in1_143 , in1_144 , in1_145 , in1_146 , in1_147 , in1_148 , in1_149 , in1_150 , in1_151 , in1_152 , in1_153 , in1_154 , in1_155 , in1_156 , in1_157 , in1_158 , in1_159 , in1_160 , in1_161 , in1_162 , in1_163 , in1_164 , in1_165 , in1_166 , in1_167 , in1_168 , in1_169 , in1_170 , in1_171 , in1_172 , in1_173 , in1_174 , in1_175 , in1_176 , in1_177 , in1_178 , in1_179 , in1_180 , in1_181 , in1_182 , in1_183 , in1_184 , in1_185 , in1_186 , in1_187 , in1_188 , in1_189 , in1_190 , in1_191 , in1_192 , in1_193 , in1_194 , in1_195 , in1_196 , in1_197 , in1_198 , in1_199 , in1_200 , in1_201 , in1_202 , in1_203 , in1_204 , in1_205 , in1_206 , in1_207 , in1_208 , in1_209 , in1_210 , in1_211 , in1_212 , in1_213 , in1_214 , in1_215 , in1_216 , in1_217 , in1_218 , in1_219 , in1_220 , in1_221 , in1_222 , in1_223 , in1_224 , in1_225 , in1_226 , in1_227 , in1_228 , in1_229 , in1_230 , in1_231 , in1_232 , in1_233 , in1_234 , in1_235 , in1_236 , in1_237 , in1_238 , in1_239 , in1_240 , in1_241 , in1_242 , in1_243 , in1_244 , in1_245 , in1_246 , in1_247 , in1_248 , in1_249 , in1_250 , in1_251 , in1_252 , in1_253 , in1_254 ,
in2_1 , in2_2 , in2_3 , in2_4 , in2_5 , in2_6 , in2_7 , in2_8 , in2_9 , in2_10 , in2_11 , in2_12 , in2_13 , in2_14 , in2_15 , in2_16 , in2_17 , in2_18 , in2_19 , in2_20 , in2_21 , in2_22 , in2_23 , in2_24 , in2_25 , in2_26 , in2_27 , in2_28 , in2_29 , in2_30 , in2_31 , in2_32 , in2_33 , in2_34 , in2_35 , in2_36 , in2_37 , in2_38 , in2_39 , in2_40 , in2_41 , in2_42 , in2_43 , in2_44 , in2_45 , in2_46 , in2_47 , in2_48 , in2_49 , in2_50 , in2_51 , in2_52 , in2_53 , in2_54 , in2_55 , in2_56 , in2_57 , in2_58 , in2_59 , in2_60 , in2_61 , in2_62 , in2_63 , in2_64 , in2_65 , in2_66 , in2_67 , in2_68 , in2_69 , in2_70 , in2_71 , in2_72 , in2_73 , in2_74 , in2_75 , in2_76 , in2_77 , in2_78 , in2_79 , in2_80 , in2_81 , in2_82 , in2_83 , in2_84 , in2_85 , in2_86 , in2_87 , in2_88 , in2_89 , in2_90 , in2_91 , in2_92 , in2_93 , in2_94 , in2_95 , in2_96 , in2_97 , in2_98 , in2_99 , in2_100 , in2_101 , in2_102 , in2_103 , in2_104 , in2_105 , in2_106 , in2_107 , in2_108 , in2_109 , in2_110 , in2_111 , in2_112 , in2_113 , in2_114 , in2_115 , in2_116 , in2_117 , in2_118 , in2_119 , in2_120 , in2_121 , in2_122 , in2_123 , in2_124 , in2_125 , in2_126 , in2_127 , in2_128 , in2_129 , in2_130 , in2_131 , in2_132 , in2_133 , in2_134 , in2_135 , in2_136 , in2_137 , in2_138 , in2_139 , in2_140 , in2_141 , in2_142 , in2_143 , in2_144 , in2_145 , in2_146 , in2_147 , in2_148 , in2_149 , in2_150 , in2_151 , in2_152 , in2_153 , in2_154 , in2_155 , in2_156 , in2_157 , in2_158 , in2_159 , in2_160 , in2_161 , in2_162 , in2_163 , in2_164 , in2_165 , in2_166 , in2_167 , in2_168 , in2_169 , in2_170 , in2_171 , in2_172 , in2_173 , in2_174 , in2_175 , in2_176 , in2_177 , in2_178 , in2_179 , in2_180 , in2_181 , in2_182 , in2_183 , in2_184 , in2_185 , in2_186 , in2_187 , in2_188 , in2_189 , in2_190 , in2_191 , in2_192 , in2_193 , in2_194 , in2_195 , in2_196 , in2_197 , in2_198 , in2_199 , in2_200 , in2_201 , in2_202 , in2_203 , in2_204 , in2_205 , in2_206 , in2_207 , in2_208 , in2_209 , in2_210 , in2_211 , in2_212 , in2_213 , in2_214 , in2_215 , in2_216 , in2_217 , in2_218 , in2_219 , in2_220 , in2_221 , in2_222 , in2_223 , in2_224 , in2_225 , in2_226 , in2_227 , in2_228 , in2_229 , in2_230 , in2_231 , in2_232 , in2_233 , in2_234 , in2_235 , in2_236 , in2_237 , in2_238 , in2_239 , in2_240 , in2_241 , in2_242 , in2_243 , in2_244 , in2_245 , in2_246 , in2_247 , in2_248 , in2_249 , in2_250 , in2_251 , in2_252 , in2_253 , in2_254 ,
out_1 , out_2 , out_3 , out_4 , out_5 , out_6 , out_7 , out_8 , out_9 , out_10 , out_11 , out_12 , out_13 , out_14 , out_15 , out_16 , out_17 , out_18 , out_19 , out_20 , out_21 , out_22 , out_23 , out_24 , out_25 , out_26 , out_27 , out_28 , out_29 , out_30 , out_31 , out_32 , out_33 , out_34 , out_35 , out_36 , out_37 , out_38 , out_39 , out_40 , out_41 , out_42 , out_43 , out_44 , out_45 , out_46 , out_47 , out_48 , out_49 , out_50 , out_51 , out_52 , out_53 , out_54 , out_55 , out_56 , out_57 , out_58 , out_59 , out_60 , out_61 , out_62 , out_63 , out_64 , out_65 , out_66 , out_67 , out_68 , out_69 , out_70 , out_71 , out_72 , out_73 , out_74 , out_75 , out_76 , out_77 , out_78 , out_79 , out_80 , out_81 , out_82 , out_83 , out_84 , out_85 , out_86 , out_87 , out_88 , out_89 , out_90 , out_91 , out_92 , out_93 , out_94 , out_95 , out_96 , out_97 , out_98 , out_99 , out_100 , out_101 , out_102 , out_103 , out_104 , out_105 , out_106 , out_107 , out_108 , out_109 , out_110 , out_111 , out_112 , out_113 , out_114 , out_115 , out_116 , out_117 , out_118 , out_119 , out_120 , out_121 , out_122 , out_123 , out_124 , out_125 , out_126 , out_127 , out_128 , out_129 , out_130 , out_131 , out_132 , out_133 , out_134 , out_135 , out_136 , out_137 , out_138 , out_139 , out_140 , out_141 , out_142 , out_143 , out_144 , out_145 , out_146 , out_147 , out_148 , out_149 , out_150 , out_151 , out_152 , out_153 , out_154 , out_155 , out_156 , out_157 , out_158 , out_159 , out_160 , out_161 , out_162 , out_163 , out_164 , out_165 , out_166 , out_167 , out_168 , out_169 , out_170 , out_171 , out_172 , out_173 , out_174 , out_175 , out_176 , out_177 , out_178 , out_179 , out_180 , out_181 , out_182 , out_183 , out_184 , out_185 , out_186 , out_187 , out_188 , out_189 , out_190 , out_191 , out_192 , out_193 , out_194 , out_195 , out_196 , out_197 , out_198 , out_199 , out_200 , out_201 , out_202 , out_203 , out_204 , out_205 , out_206 , out_207 , out_208 , out_209 , out_210 , out_211 , out_212 , out_213 , out_214 , out_215 , out_216 , out_217 , out_218 , out_219 , out_220 , out_221 , out_222 , out_223 , out_224 , out_225 , out_226 , out_227 , out_228 , out_229 , out_230 , out_231 , out_232 , out_233 , out_234 , out_235 , out_236 , out_237 , out_238 , out_239 , out_240 , out_241 , out_242 , out_243 , out_244 , out_245 , out_246 , out_247 , out_248 , out_249 , out_250 , out_251 , out_252 , out_253 , out_254 
);

input in1_1 , in1_2 , in1_3 , in1_4 , in1_5 , in1_6 , in1_7 , in1_8 , in1_9 , in1_10 , in1_11 , in1_12 , in1_13 , in1_14 , in1_15 , in1_16 , in1_17 , in1_18 , in1_19 , in1_20 , in1_21 , in1_22 , in1_23 , in1_24 , in1_25 , in1_26 , in1_27 , in1_28 , in1_29 , in1_30 , in1_31 , in1_32 , in1_33 , in1_34 , in1_35 , in1_36 , in1_37 , in1_38 , in1_39 , in1_40 , in1_41 , in1_42 , in1_43 , in1_44 , in1_45 , in1_46 , in1_47 , in1_48 , in1_49 , in1_50 , in1_51 , in1_52 , in1_53 , in1_54 , in1_55 , in1_56 , in1_57 , in1_58 , in1_59 , in1_60 , in1_61 , in1_62 , in1_63 , in1_64 , in1_65 , in1_66 , in1_67 , in1_68 , in1_69 , in1_70 , in1_71 , in1_72 , in1_73 , in1_74 , in1_75 , in1_76 , in1_77 , in1_78 , in1_79 , in1_80 , in1_81 , in1_82 , in1_83 , in1_84 , in1_85 , in1_86 , in1_87 , in1_88 , in1_89 , in1_90 , in1_91 , in1_92 , in1_93 , in1_94 , in1_95 , in1_96 , in1_97 , in1_98 , in1_99 , in1_100 , in1_101 , in1_102 , in1_103 , in1_104 , in1_105 , in1_106 , in1_107 , in1_108 , in1_109 , in1_110 , in1_111 , in1_112 , in1_113 , in1_114 , in1_115 , in1_116 , in1_117 , in1_118 , in1_119 , in1_120 , in1_121 , in1_122 , in1_123 , in1_124 , in1_125 , in1_126 , in1_127 , in1_128 , in1_129 , in1_130 , in1_131 , in1_132 , in1_133 , in1_134 , in1_135 , in1_136 , in1_137 , in1_138 , in1_139 , in1_140 , in1_141 , in1_142 , in1_143 , in1_144 , in1_145 , in1_146 , in1_147 , in1_148 , in1_149 , in1_150 , in1_151 , in1_152 , in1_153 , in1_154 , in1_155 , in1_156 , in1_157 , in1_158 , in1_159 , in1_160 , in1_161 , in1_162 , in1_163 , in1_164 , in1_165 , in1_166 , in1_167 , in1_168 , in1_169 , in1_170 , in1_171 , in1_172 , in1_173 , in1_174 , in1_175 , in1_176 , in1_177 , in1_178 , in1_179 , in1_180 , in1_181 , in1_182 , in1_183 , in1_184 , in1_185 , in1_186 , in1_187 , in1_188 , in1_189 , in1_190 , in1_191 , in1_192 , in1_193 , in1_194 , in1_195 , in1_196 , in1_197 , in1_198 , in1_199 , in1_200 , in1_201 , in1_202 , in1_203 , in1_204 , in1_205 , in1_206 , in1_207 , in1_208 , in1_209 , in1_210 , in1_211 , in1_212 , in1_213 , in1_214 , in1_215 , in1_216 , in1_217 , in1_218 , in1_219 , in1_220 , in1_221 , in1_222 , in1_223 , in1_224 , in1_225 , in1_226 , in1_227 , in1_228 , in1_229 , in1_230 , in1_231 , in1_232 , in1_233 , in1_234 , in1_235 , in1_236 , in1_237 , in1_238 , in1_239 , in1_240 , in1_241 , in1_242 , in1_243 , in1_244 , in1_245 , in1_246 , in1_247 , in1_248 , in1_249 , in1_250 , in1_251 , in1_252 , in1_253 , in1_254 ;
input in2_1 , in2_2 , in2_3 , in2_4 , in2_5 , in2_6 , in2_7 , in2_8 , in2_9 , in2_10 , in2_11 , in2_12 , in2_13 , in2_14 , in2_15 , in2_16 , in2_17 , in2_18 , in2_19 , in2_20 , in2_21 , in2_22 , in2_23 , in2_24 , in2_25 , in2_26 , in2_27 , in2_28 , in2_29 , in2_30 , in2_31 , in2_32 , in2_33 , in2_34 , in2_35 , in2_36 , in2_37 , in2_38 , in2_39 , in2_40 , in2_41 , in2_42 , in2_43 , in2_44 , in2_45 , in2_46 , in2_47 , in2_48 , in2_49 , in2_50 , in2_51 , in2_52 , in2_53 , in2_54 , in2_55 , in2_56 , in2_57 , in2_58 , in2_59 , in2_60 , in2_61 , in2_62 , in2_63 , in2_64 , in2_65 , in2_66 , in2_67 , in2_68 , in2_69 , in2_70 , in2_71 , in2_72 , in2_73 , in2_74 , in2_75 , in2_76 , in2_77 , in2_78 , in2_79 , in2_80 , in2_81 , in2_82 , in2_83 , in2_84 , in2_85 , in2_86 , in2_87 , in2_88 , in2_89 , in2_90 , in2_91 , in2_92 , in2_93 , in2_94 , in2_95 , in2_96 , in2_97 , in2_98 , in2_99 , in2_100 , in2_101 , in2_102 , in2_103 , in2_104 , in2_105 , in2_106 , in2_107 , in2_108 , in2_109 , in2_110 , in2_111 , in2_112 , in2_113 , in2_114 , in2_115 , in2_116 , in2_117 , in2_118 , in2_119 , in2_120 , in2_121 , in2_122 , in2_123 , in2_124 , in2_125 , in2_126 , in2_127 , in2_128 , in2_129 , in2_130 , in2_131 , in2_132 , in2_133 , in2_134 , in2_135 , in2_136 , in2_137 , in2_138 , in2_139 , in2_140 , in2_141 , in2_142 , in2_143 , in2_144 , in2_145 , in2_146 , in2_147 , in2_148 , in2_149 , in2_150 , in2_151 , in2_152 , in2_153 , in2_154 , in2_155 , in2_156 , in2_157 , in2_158 , in2_159 , in2_160 , in2_161 , in2_162 , in2_163 , in2_164 , in2_165 , in2_166 , in2_167 , in2_168 , in2_169 , in2_170 , in2_171 , in2_172 , in2_173 , in2_174 , in2_175 , in2_176 , in2_177 , in2_178 , in2_179 , in2_180 , in2_181 , in2_182 , in2_183 , in2_184 , in2_185 , in2_186 , in2_187 , in2_188 , in2_189 , in2_190 , in2_191 , in2_192 , in2_193 , in2_194 , in2_195 , in2_196 , in2_197 , in2_198 , in2_199 , in2_200 , in2_201 , in2_202 , in2_203 , in2_204 , in2_205 , in2_206 , in2_207 , in2_208 , in2_209 , in2_210 , in2_211 , in2_212 , in2_213 , in2_214 , in2_215 , in2_216 , in2_217 , in2_218 , in2_219 , in2_220 , in2_221 , in2_222 , in2_223 , in2_224 , in2_225 , in2_226 , in2_227 , in2_228 , in2_229 , in2_230 , in2_231 , in2_232 , in2_233 , in2_234 , in2_235 , in2_236 , in2_237 , in2_238 , in2_239 , in2_240 , in2_241 , in2_242 , in2_243 , in2_244 , in2_245 , in2_246 , in2_247 , in2_248 , in2_249 , in2_250 , in2_251 , in2_252 , in2_253 , in2_254 ;

output out_1 , out_2 , out_3 , out_4 , out_5 , out_6 , out_7 , out_8 , out_9 , out_10 , out_11 , out_12 , out_13 , out_14 , out_15 , out_16 , out_17 , out_18 , out_19 , out_20 , out_21 , out_22 , out_23 , out_24 , out_25 , out_26 , out_27 , out_28 , out_29 , out_30 , out_31 , out_32 , out_33 , out_34 , out_35 , out_36 , out_37 , out_38 , out_39 , out_40 , out_41 , out_42 , out_43 , out_44 , out_45 , out_46 , out_47 , out_48 , out_49 , out_50 , out_51 , out_52 , out_53 , out_54 , out_55 , out_56 , out_57 , out_58 , out_59 , out_60 , out_61 , out_62 , out_63 , out_64 , out_65 , out_66 , out_67 , out_68 , out_69 , out_70 , out_71 , out_72 , out_73 , out_74 , out_75 , out_76 , out_77 , out_78 , out_79 , out_80 , out_81 , out_82 , out_83 , out_84 , out_85 , out_86 , out_87 , out_88 , out_89 , out_90 , out_91 , out_92 , out_93 , out_94 , out_95 , out_96 , out_97 , out_98 , out_99 , out_100 , out_101 , out_102 , out_103 , out_104 , out_105 , out_106 , out_107 , out_108 , out_109 , out_110 , out_111 , out_112 , out_113 , out_114 , out_115 , out_116 , out_117 , out_118 , out_119 , out_120 , out_121 , out_122 , out_123 , out_124 , out_125 , out_126 , out_127 , out_128 , out_129 , out_130 , out_131 , out_132 , out_133 , out_134 , out_135 , out_136 , out_137 , out_138 , out_139 , out_140 , out_141 , out_142 , out_143 , out_144 , out_145 , out_146 , out_147 , out_148 , out_149 , out_150 , out_151 , out_152 , out_153 , out_154 , out_155 , out_156 , out_157 , out_158 , out_159 , out_160 , out_161 , out_162 , out_163 , out_164 , out_165 , out_166 , out_167 , out_168 , out_169 , out_170 , out_171 , out_172 , out_173 , out_174 , out_175 , out_176 , out_177 , out_178 , out_179 , out_180 , out_181 , out_182 , out_183 , out_184 , out_185 , out_186 , out_187 , out_188 , out_189 , out_190 , out_191 , out_192 , out_193 , out_194 , out_195 , out_196 , out_197 , out_198 , out_199 , out_200 , out_201 , out_202 , out_203 , out_204 , out_205 , out_206 , out_207 , out_208 , out_209 , out_210 , out_211 , out_212 , out_213 , out_214 , out_215 , out_216 , out_217 , out_218 , out_219 , out_220 , out_221 , out_222 , out_223 , out_224 , out_225 , out_226 , out_227 , out_228 , out_229 , out_230 , out_231 , out_232 , out_233 , out_234 , out_235 , out_236 , out_237 , out_238 , out_239 , out_240 , out_241 , out_242 , out_243 , out_244 , out_245 , out_246 , out_247 , out_248 , out_249 , out_250 , out_251 , out_252 , out_253 , out_254 ;


assign out_1 = in1_1 ^ in2_1 ; 
assign out_2 = in1_2 ^ in2_2 ; 
assign out_3 = in1_3 ^ in2_3 ; 
assign out_4 = in1_4 ^ in2_4 ; 
assign out_5 = in1_5 ^ in2_5 ; 
assign out_6 = in1_6 ^ in2_6 ; 
assign out_7 = in1_7 ^ in2_7 ; 
assign out_8 = in1_8 ^ in2_8 ; 
assign out_9 = in1_9 ^ in2_9 ; 
assign out_10 = in1_10 ^ in2_10 ; 
assign out_11 = in1_11 ^ in2_11 ; 
assign out_12 = in1_12 ^ in2_12 ; 
assign out_13 = in1_13 ^ in2_13 ; 
assign out_14 = in1_14 ^ in2_14 ; 
assign out_15 = in1_15 ^ in2_15 ; 
assign out_16 = in1_16 ^ in2_16 ; 
assign out_17 = in1_17 ^ in2_17 ; 
assign out_18 = in1_18 ^ in2_18 ; 
assign out_19 = in1_19 ^ in2_19 ; 
assign out_20 = in1_20 ^ in2_20 ; 
assign out_21 = in1_21 ^ in2_21 ; 
assign out_22 = in1_22 ^ in2_22 ; 
assign out_23 = in1_23 ^ in2_23 ; 
assign out_24 = in1_24 ^ in2_24 ; 
assign out_25 = in1_25 ^ in2_25 ; 
assign out_26 = in1_26 ^ in2_26 ; 
assign out_27 = in1_27 ^ in2_27 ; 
assign out_28 = in1_28 ^ in2_28 ; 
assign out_29 = in1_29 ^ in2_29 ; 
assign out_30 = in1_30 ^ in2_30 ; 
assign out_31 = in1_31 ^ in2_31 ; 
assign out_32 = in1_32 ^ in2_32 ; 
assign out_33 = in1_33 ^ in2_33 ; 
assign out_34 = in1_34 ^ in2_34 ; 
assign out_35 = in1_35 ^ in2_35 ; 
assign out_36 = in1_36 ^ in2_36 ; 
assign out_37 = in1_37 ^ in2_37 ; 
assign out_38 = in1_38 ^ in2_38 ; 
assign out_39 = in1_39 ^ in2_39 ; 
assign out_40 = in1_40 ^ in2_40 ; 
assign out_41 = in1_41 ^ in2_41 ; 
assign out_42 = in1_42 ^ in2_42 ; 
assign out_43 = in1_43 ^ in2_43 ; 
assign out_44 = in1_44 ^ in2_44 ; 
assign out_45 = in1_45 ^ in2_45 ; 
assign out_46 = in1_46 ^ in2_46 ; 
assign out_47 = in1_47 ^ in2_47 ; 
assign out_48 = in1_48 ^ in2_48 ; 
assign out_49 = in1_49 ^ in2_49 ; 
assign out_50 = in1_50 ^ in2_50 ; 
assign out_51 = in1_51 ^ in2_51 ; 
assign out_52 = in1_52 ^ in2_52 ; 
assign out_53 = in1_53 ^ in2_53 ; 
assign out_54 = in1_54 ^ in2_54 ; 
assign out_55 = in1_55 ^ in2_55 ; 
assign out_56 = in1_56 ^ in2_56 ; 
assign out_57 = in1_57 ^ in2_57 ; 
assign out_58 = in1_58 ^ in2_58 ; 
assign out_59 = in1_59 ^ in2_59 ; 
assign out_60 = in1_60 ^ in2_60 ; 
assign out_61 = in1_61 ^ in2_61 ; 
assign out_62 = in1_62 ^ in2_62 ; 
assign out_63 = in1_63 ^ in2_63 ; 
assign out_64 = in1_64 ^ in2_64 ; 
assign out_65 = in1_65 ^ in2_65 ; 
assign out_66 = in1_66 ^ in2_66 ; 
assign out_67 = in1_67 ^ in2_67 ; 
assign out_68 = in1_68 ^ in2_68 ; 
assign out_69 = in1_69 ^ in2_69 ; 
assign out_70 = in1_70 ^ in2_70 ; 
assign out_71 = in1_71 ^ in2_71 ; 
assign out_72 = in1_72 ^ in2_72 ; 
assign out_73 = in1_73 ^ in2_73 ; 
assign out_74 = in1_74 ^ in2_74 ; 
assign out_75 = in1_75 ^ in2_75 ; 
assign out_76 = in1_76 ^ in2_76 ; 
assign out_77 = in1_77 ^ in2_77 ; 
assign out_78 = in1_78 ^ in2_78 ; 
assign out_79 = in1_79 ^ in2_79 ; 
assign out_80 = in1_80 ^ in2_80 ; 
assign out_81 = in1_81 ^ in2_81 ; 
assign out_82 = in1_82 ^ in2_82 ; 
assign out_83 = in1_83 ^ in2_83 ; 
assign out_84 = in1_84 ^ in2_84 ; 
assign out_85 = in1_85 ^ in2_85 ; 
assign out_86 = in1_86 ^ in2_86 ; 
assign out_87 = in1_87 ^ in2_87 ; 
assign out_88 = in1_88 ^ in2_88 ; 
assign out_89 = in1_89 ^ in2_89 ; 
assign out_90 = in1_90 ^ in2_90 ; 
assign out_91 = in1_91 ^ in2_91 ; 
assign out_92 = in1_92 ^ in2_92 ; 
assign out_93 = in1_93 ^ in2_93 ; 
assign out_94 = in1_94 ^ in2_94 ; 
assign out_95 = in1_95 ^ in2_95 ; 
assign out_96 = in1_96 ^ in2_96 ; 
assign out_97 = in1_97 ^ in2_97 ; 
assign out_98 = in1_98 ^ in2_98 ; 
assign out_99 = in1_99 ^ in2_99 ; 
assign out_100 = in1_100 ^ in2_100 ; 
assign out_101 = in1_101 ^ in2_101 ; 
assign out_102 = in1_102 ^ in2_102 ; 
assign out_103 = in1_103 ^ in2_103 ; 
assign out_104 = in1_104 ^ in2_104 ; 
assign out_105 = in1_105 ^ in2_105 ; 
assign out_106 = in1_106 ^ in2_106 ; 
assign out_107 = in1_107 ^ in2_107 ; 
assign out_108 = in1_108 ^ in2_108 ; 
assign out_109 = in1_109 ^ in2_109 ; 
assign out_110 = in1_110 ^ in2_110 ; 
assign out_111 = in1_111 ^ in2_111 ; 
assign out_112 = in1_112 ^ in2_112 ; 
assign out_113 = in1_113 ^ in2_113 ; 
assign out_114 = in1_114 ^ in2_114 ; 
assign out_115 = in1_115 ^ in2_115 ; 
assign out_116 = in1_116 ^ in2_116 ; 
assign out_117 = in1_117 ^ in2_117 ; 
assign out_118 = in1_118 ^ in2_118 ; 
assign out_119 = in1_119 ^ in2_119 ; 
assign out_120 = in1_120 ^ in2_120 ; 
assign out_121 = in1_121 ^ in2_121 ; 
assign out_122 = in1_122 ^ in2_122 ; 
assign out_123 = in1_123 ^ in2_123 ; 
assign out_124 = in1_124 ^ in2_124 ; 
assign out_125 = in1_125 ^ in2_125 ; 
assign out_126 = in1_126 ^ in2_126 ; 
assign out_127 = in1_127 ^ in2_127 ; 
assign out_128 = in1_128 ^ in2_128 ; 
assign out_129 = in1_129 ^ in2_129 ; 
assign out_130 = in1_130 ^ in2_130 ; 
assign out_131 = in1_131 ^ in2_131 ; 
assign out_132 = in1_132 ^ in2_132 ; 
assign out_133 = in1_133 ^ in2_133 ; 
assign out_134 = in1_134 ^ in2_134 ; 
assign out_135 = in1_135 ^ in2_135 ; 
assign out_136 = in1_136 ^ in2_136 ; 
assign out_137 = in1_137 ^ in2_137 ; 
assign out_138 = in1_138 ^ in2_138 ; 
assign out_139 = in1_139 ^ in2_139 ; 
assign out_140 = in1_140 ^ in2_140 ; 
assign out_141 = in1_141 ^ in2_141 ; 
assign out_142 = in1_142 ^ in2_142 ; 
assign out_143 = in1_143 ^ in2_143 ; 
assign out_144 = in1_144 ^ in2_144 ; 
assign out_145 = in1_145 ^ in2_145 ; 
assign out_146 = in1_146 ^ in2_146 ; 
assign out_147 = in1_147 ^ in2_147 ; 
assign out_148 = in1_148 ^ in2_148 ; 
assign out_149 = in1_149 ^ in2_149 ; 
assign out_150 = in1_150 ^ in2_150 ; 
assign out_151 = in1_151 ^ in2_151 ; 
assign out_152 = in1_152 ^ in2_152 ; 
assign out_153 = in1_153 ^ in2_153 ; 
assign out_154 = in1_154 ^ in2_154 ; 
assign out_155 = in1_155 ^ in2_155 ; 
assign out_156 = in1_156 ^ in2_156 ; 
assign out_157 = in1_157 ^ in2_157 ; 
assign out_158 = in1_158 ^ in2_158 ; 
assign out_159 = in1_159 ^ in2_159 ; 
assign out_160 = in1_160 ^ in2_160 ; 
assign out_161 = in1_161 ^ in2_161 ; 
assign out_162 = in1_162 ^ in2_162 ; 
assign out_163 = in1_163 ^ in2_163 ; 
assign out_164 = in1_164 ^ in2_164 ; 
assign out_165 = in1_165 ^ in2_165 ; 
assign out_166 = in1_166 ^ in2_166 ; 
assign out_167 = in1_167 ^ in2_167 ; 
assign out_168 = in1_168 ^ in2_168 ; 
assign out_169 = in1_169 ^ in2_169 ; 
assign out_170 = in1_170 ^ in2_170 ; 
assign out_171 = in1_171 ^ in2_171 ; 
assign out_172 = in1_172 ^ in2_172 ; 
assign out_173 = in1_173 ^ in2_173 ; 
assign out_174 = in1_174 ^ in2_174 ; 
assign out_175 = in1_175 ^ in2_175 ; 
assign out_176 = in1_176 ^ in2_176 ; 
assign out_177 = in1_177 ^ in2_177 ; 
assign out_178 = in1_178 ^ in2_178 ; 
assign out_179 = in1_179 ^ in2_179 ; 
assign out_180 = in1_180 ^ in2_180 ; 
assign out_181 = in1_181 ^ in2_181 ; 
assign out_182 = in1_182 ^ in2_182 ; 
assign out_183 = in1_183 ^ in2_183 ; 
assign out_184 = in1_184 ^ in2_184 ; 
assign out_185 = in1_185 ^ in2_185 ; 
assign out_186 = in1_186 ^ in2_186 ; 
assign out_187 = in1_187 ^ in2_187 ; 
assign out_188 = in1_188 ^ in2_188 ; 
assign out_189 = in1_189 ^ in2_189 ; 
assign out_190 = in1_190 ^ in2_190 ; 
assign out_191 = in1_191 ^ in2_191 ; 
assign out_192 = in1_192 ^ in2_192 ; 
assign out_193 = in1_193 ^ in2_193 ; 
assign out_194 = in1_194 ^ in2_194 ; 
assign out_195 = in1_195 ^ in2_195 ; 
assign out_196 = in1_196 ^ in2_196 ; 
assign out_197 = in1_197 ^ in2_197 ; 
assign out_198 = in1_198 ^ in2_198 ; 
assign out_199 = in1_199 ^ in2_199 ; 
assign out_200 = in1_200 ^ in2_200 ; 
assign out_201 = in1_201 ^ in2_201 ; 
assign out_202 = in1_202 ^ in2_202 ; 
assign out_203 = in1_203 ^ in2_203 ; 
assign out_204 = in1_204 ^ in2_204 ; 
assign out_205 = in1_205 ^ in2_205 ; 
assign out_206 = in1_206 ^ in2_206 ; 
assign out_207 = in1_207 ^ in2_207 ; 
assign out_208 = in1_208 ^ in2_208 ; 
assign out_209 = in1_209 ^ in2_209 ; 
assign out_210 = in1_210 ^ in2_210 ; 
assign out_211 = in1_211 ^ in2_211 ; 
assign out_212 = in1_212 ^ in2_212 ; 
assign out_213 = in1_213 ^ in2_213 ; 
assign out_214 = in1_214 ^ in2_214 ; 
assign out_215 = in1_215 ^ in2_215 ; 
assign out_216 = in1_216 ^ in2_216 ; 
assign out_217 = in1_217 ^ in2_217 ; 
assign out_218 = in1_218 ^ in2_218 ; 
assign out_219 = in1_219 ^ in2_219 ; 
assign out_220 = in1_220 ^ in2_220 ; 
assign out_221 = in1_221 ^ in2_221 ; 
assign out_222 = in1_222 ^ in2_222 ; 
assign out_223 = in1_223 ^ in2_223 ; 
assign out_224 = in1_224 ^ in2_224 ; 
assign out_225 = in1_225 ^ in2_225 ; 
assign out_226 = in1_226 ^ in2_226 ; 
assign out_227 = in1_227 ^ in2_227 ; 
assign out_228 = in1_228 ^ in2_228 ; 
assign out_229 = in1_229 ^ in2_229 ; 
assign out_230 = in1_230 ^ in2_230 ; 
assign out_231 = in1_231 ^ in2_231 ; 
assign out_232 = in1_232 ^ in2_232 ; 
assign out_233 = in1_233 ^ in2_233 ; 
assign out_234 = in1_234 ^ in2_234 ; 
assign out_235 = in1_235 ^ in2_235 ; 
assign out_236 = in1_236 ^ in2_236 ; 
assign out_237 = in1_237 ^ in2_237 ; 
assign out_238 = in1_238 ^ in2_238 ; 
assign out_239 = in1_239 ^ in2_239 ; 
assign out_240 = in1_240 ^ in2_240 ; 
assign out_241 = in1_241 ^ in2_241 ; 
assign out_242 = in1_242 ^ in2_242 ; 
assign out_243 = in1_243 ^ in2_243 ; 
assign out_244 = in1_244 ^ in2_244 ; 
assign out_245 = in1_245 ^ in2_245 ; 
assign out_246 = in1_246 ^ in2_246 ; 
assign out_247 = in1_247 ^ in2_247 ; 
assign out_248 = in1_248 ^ in2_248 ; 
assign out_249 = in1_249 ^ in2_249 ; 
assign out_250 = in1_250 ^ in2_250 ; 
assign out_251 = in1_251 ^ in2_251 ; 
assign out_252 = in1_252 ^ in2_252 ; 
assign out_253 = in1_253 ^ in2_253 ; 
assign out_254 = in1_254 ^ in2_254 ; 

endmodule