`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 02/22/2025
// Design Name: sum_of_second_module_outputs
// Module Name: sum_of_second_module_outputs
// Description: This module calculates the sum of various shares from the second module.
//              It computes sums based on specific equations related to cross-module terms.
// Dependencies: None
// Revision: 0.01 - Initial version
//////////////////////////////////////////////////////////////////////////////////

module sum_of_second_module_outputs (
    output_x4_share ,  output_x5_share ,  output_x6_share ,  output_x7_share ,  output_x4x5_share ,  output_x4x6_share ,  output_x4x7_share ,  output_x5x6_share ,  output_x5x7_share ,  output_x6x7_share ,  output_x4x5x6_share ,  output_x4x5x7_share ,  output_x4x6x7_share ,  output_x5x6x7_share ,  output_x4x5x6x7_share,
output_sum_secondmodule_equation_num_0_index_0_share, output_sum_secondmodule_equation_num_0_index_1_share, output_sum_secondmodule_equation_num_0_index_2_share, output_sum_secondmodule_equation_num_0_index_3_share, output_sum_secondmodule_equation_num_0_index_4_share, output_sum_secondmodule_equation_num_0_index_5_share, output_sum_secondmodule_equation_num_0_index_6_share, output_sum_secondmodule_equation_num_0_index_7_share, output_sum_secondmodule_equation_num_0_index_8_share, output_sum_secondmodule_equation_num_0_index_9_share, output_sum_secondmodule_equation_num_0_index_10_share, output_sum_secondmodule_equation_num_0_index_11_share, output_sum_secondmodule_equation_num_0_index_12_share, output_sum_secondmodule_equation_num_0_index_13_share, output_sum_secondmodule_equation_num_0_index_14_share,
output_sum_secondmodule_equation_num_1_index_0_share, output_sum_secondmodule_equation_num_1_index_1_share, output_sum_secondmodule_equation_num_1_index_2_share, output_sum_secondmodule_equation_num_1_index_3_share, output_sum_secondmodule_equation_num_1_index_4_share, output_sum_secondmodule_equation_num_1_index_5_share, output_sum_secondmodule_equation_num_1_index_6_share, output_sum_secondmodule_equation_num_1_index_7_share, output_sum_secondmodule_equation_num_1_index_8_share, output_sum_secondmodule_equation_num_1_index_9_share, output_sum_secondmodule_equation_num_1_index_10_share, output_sum_secondmodule_equation_num_1_index_11_share, output_sum_secondmodule_equation_num_1_index_12_share, output_sum_secondmodule_equation_num_1_index_13_share, output_sum_secondmodule_equation_num_1_index_14_share,
output_sum_secondmodule_equation_num_2_index_0_share, output_sum_secondmodule_equation_num_2_index_1_share, output_sum_secondmodule_equation_num_2_index_2_share, output_sum_secondmodule_equation_num_2_index_3_share, output_sum_secondmodule_equation_num_2_index_4_share, output_sum_secondmodule_equation_num_2_index_5_share, output_sum_secondmodule_equation_num_2_index_6_share, output_sum_secondmodule_equation_num_2_index_7_share, output_sum_secondmodule_equation_num_2_index_8_share, output_sum_secondmodule_equation_num_2_index_9_share, output_sum_secondmodule_equation_num_2_index_10_share, output_sum_secondmodule_equation_num_2_index_11_share, output_sum_secondmodule_equation_num_2_index_12_share, output_sum_secondmodule_equation_num_2_index_13_share, output_sum_secondmodule_equation_num_2_index_14_share,
output_sum_secondmodule_equation_num_3_index_0_share, output_sum_secondmodule_equation_num_3_index_1_share, output_sum_secondmodule_equation_num_3_index_2_share, output_sum_secondmodule_equation_num_3_index_3_share, output_sum_secondmodule_equation_num_3_index_4_share, output_sum_secondmodule_equation_num_3_index_5_share, output_sum_secondmodule_equation_num_3_index_6_share, output_sum_secondmodule_equation_num_3_index_7_share, output_sum_secondmodule_equation_num_3_index_8_share, output_sum_secondmodule_equation_num_3_index_9_share, output_sum_secondmodule_equation_num_3_index_10_share, output_sum_secondmodule_equation_num_3_index_11_share, output_sum_secondmodule_equation_num_3_index_12_share, output_sum_secondmodule_equation_num_3_index_13_share, output_sum_secondmodule_equation_num_3_index_14_share,
output_sum_secondmodule_equation_num_4_index_0_share, output_sum_secondmodule_equation_num_4_index_1_share, output_sum_secondmodule_equation_num_4_index_2_share, output_sum_secondmodule_equation_num_4_index_3_share, output_sum_secondmodule_equation_num_4_index_4_share, output_sum_secondmodule_equation_num_4_index_5_share, output_sum_secondmodule_equation_num_4_index_6_share, output_sum_secondmodule_equation_num_4_index_7_share, output_sum_secondmodule_equation_num_4_index_8_share, output_sum_secondmodule_equation_num_4_index_9_share, output_sum_secondmodule_equation_num_4_index_10_share, output_sum_secondmodule_equation_num_4_index_11_share, output_sum_secondmodule_equation_num_4_index_12_share, output_sum_secondmodule_equation_num_4_index_13_share, output_sum_secondmodule_equation_num_4_index_14_share,
output_sum_secondmodule_equation_num_5_index_0_share, output_sum_secondmodule_equation_num_5_index_1_share, output_sum_secondmodule_equation_num_5_index_2_share, output_sum_secondmodule_equation_num_5_index_3_share, output_sum_secondmodule_equation_num_5_index_4_share, output_sum_secondmodule_equation_num_5_index_5_share, output_sum_secondmodule_equation_num_5_index_6_share, output_sum_secondmodule_equation_num_5_index_7_share, output_sum_secondmodule_equation_num_5_index_8_share, output_sum_secondmodule_equation_num_5_index_9_share, output_sum_secondmodule_equation_num_5_index_10_share, output_sum_secondmodule_equation_num_5_index_11_share, output_sum_secondmodule_equation_num_5_index_12_share, output_sum_secondmodule_equation_num_5_index_13_share, output_sum_secondmodule_equation_num_5_index_14_share,
output_sum_secondmodule_equation_num_6_index_0_share, output_sum_secondmodule_equation_num_6_index_1_share, output_sum_secondmodule_equation_num_6_index_2_share, output_sum_secondmodule_equation_num_6_index_3_share, output_sum_secondmodule_equation_num_6_index_4_share, output_sum_secondmodule_equation_num_6_index_5_share, output_sum_secondmodule_equation_num_6_index_6_share, output_sum_secondmodule_equation_num_6_index_7_share, output_sum_secondmodule_equation_num_6_index_8_share, output_sum_secondmodule_equation_num_6_index_9_share, output_sum_secondmodule_equation_num_6_index_10_share, output_sum_secondmodule_equation_num_6_index_11_share, output_sum_secondmodule_equation_num_6_index_12_share, output_sum_secondmodule_equation_num_6_index_13_share, output_sum_secondmodule_equation_num_6_index_14_share,
output_sum_secondmodule_equation_num_7_index_0_share, output_sum_secondmodule_equation_num_7_index_1_share, output_sum_secondmodule_equation_num_7_index_2_share, output_sum_secondmodule_equation_num_7_index_3_share, output_sum_secondmodule_equation_num_7_index_4_share, output_sum_secondmodule_equation_num_7_index_5_share, output_sum_secondmodule_equation_num_7_index_6_share, output_sum_secondmodule_equation_num_7_index_7_share, output_sum_secondmodule_equation_num_7_index_8_share, output_sum_secondmodule_equation_num_7_index_9_share, output_sum_secondmodule_equation_num_7_index_10_share, output_sum_secondmodule_equation_num_7_index_11_share, output_sum_secondmodule_equation_num_7_index_12_share, output_sum_secondmodule_equation_num_7_index_13_share, output_sum_secondmodule_equation_num_7_index_14_share

);

input  output_x4_share ,  output_x5_share ,  output_x6_share ,  output_x7_share ,  output_x4x5_share ,  output_x4x6_share ,  output_x4x7_share ,  output_x5x6_share ,  output_x5x7_share ,  output_x6x7_share ,  output_x4x5x6_share ,  output_x4x5x7_share ,  output_x4x6x7_share ,  output_x5x6x7_share ,  output_x4x5x6x7_share ;
output output_sum_secondmodule_equation_num_0_index_0_share, output_sum_secondmodule_equation_num_0_index_1_share, output_sum_secondmodule_equation_num_0_index_2_share, output_sum_secondmodule_equation_num_0_index_3_share, output_sum_secondmodule_equation_num_0_index_4_share, output_sum_secondmodule_equation_num_0_index_5_share, output_sum_secondmodule_equation_num_0_index_6_share, output_sum_secondmodule_equation_num_0_index_7_share, output_sum_secondmodule_equation_num_0_index_8_share, output_sum_secondmodule_equation_num_0_index_9_share, output_sum_secondmodule_equation_num_0_index_10_share, output_sum_secondmodule_equation_num_0_index_11_share, output_sum_secondmodule_equation_num_0_index_12_share, output_sum_secondmodule_equation_num_0_index_13_share, output_sum_secondmodule_equation_num_0_index_14_share;
output output_sum_secondmodule_equation_num_1_index_0_share, output_sum_secondmodule_equation_num_1_index_1_share, output_sum_secondmodule_equation_num_1_index_2_share, output_sum_secondmodule_equation_num_1_index_3_share, output_sum_secondmodule_equation_num_1_index_4_share, output_sum_secondmodule_equation_num_1_index_5_share, output_sum_secondmodule_equation_num_1_index_6_share, output_sum_secondmodule_equation_num_1_index_7_share, output_sum_secondmodule_equation_num_1_index_8_share, output_sum_secondmodule_equation_num_1_index_9_share, output_sum_secondmodule_equation_num_1_index_10_share, output_sum_secondmodule_equation_num_1_index_11_share, output_sum_secondmodule_equation_num_1_index_12_share, output_sum_secondmodule_equation_num_1_index_13_share, output_sum_secondmodule_equation_num_1_index_14_share;
output output_sum_secondmodule_equation_num_2_index_0_share, output_sum_secondmodule_equation_num_2_index_1_share, output_sum_secondmodule_equation_num_2_index_2_share, output_sum_secondmodule_equation_num_2_index_3_share, output_sum_secondmodule_equation_num_2_index_4_share, output_sum_secondmodule_equation_num_2_index_5_share, output_sum_secondmodule_equation_num_2_index_6_share, output_sum_secondmodule_equation_num_2_index_7_share, output_sum_secondmodule_equation_num_2_index_8_share, output_sum_secondmodule_equation_num_2_index_9_share, output_sum_secondmodule_equation_num_2_index_10_share, output_sum_secondmodule_equation_num_2_index_11_share, output_sum_secondmodule_equation_num_2_index_12_share, output_sum_secondmodule_equation_num_2_index_13_share, output_sum_secondmodule_equation_num_2_index_14_share;
output output_sum_secondmodule_equation_num_3_index_0_share, output_sum_secondmodule_equation_num_3_index_1_share, output_sum_secondmodule_equation_num_3_index_2_share, output_sum_secondmodule_equation_num_3_index_3_share, output_sum_secondmodule_equation_num_3_index_4_share, output_sum_secondmodule_equation_num_3_index_5_share, output_sum_secondmodule_equation_num_3_index_6_share, output_sum_secondmodule_equation_num_3_index_7_share, output_sum_secondmodule_equation_num_3_index_8_share, output_sum_secondmodule_equation_num_3_index_9_share, output_sum_secondmodule_equation_num_3_index_10_share, output_sum_secondmodule_equation_num_3_index_11_share, output_sum_secondmodule_equation_num_3_index_12_share, output_sum_secondmodule_equation_num_3_index_13_share, output_sum_secondmodule_equation_num_3_index_14_share;
output output_sum_secondmodule_equation_num_4_index_0_share, output_sum_secondmodule_equation_num_4_index_1_share, output_sum_secondmodule_equation_num_4_index_2_share, output_sum_secondmodule_equation_num_4_index_3_share, output_sum_secondmodule_equation_num_4_index_4_share, output_sum_secondmodule_equation_num_4_index_5_share, output_sum_secondmodule_equation_num_4_index_6_share, output_sum_secondmodule_equation_num_4_index_7_share, output_sum_secondmodule_equation_num_4_index_8_share, output_sum_secondmodule_equation_num_4_index_9_share, output_sum_secondmodule_equation_num_4_index_10_share, output_sum_secondmodule_equation_num_4_index_11_share, output_sum_secondmodule_equation_num_4_index_12_share, output_sum_secondmodule_equation_num_4_index_13_share, output_sum_secondmodule_equation_num_4_index_14_share;
output output_sum_secondmodule_equation_num_5_index_0_share, output_sum_secondmodule_equation_num_5_index_1_share, output_sum_secondmodule_equation_num_5_index_2_share, output_sum_secondmodule_equation_num_5_index_3_share, output_sum_secondmodule_equation_num_5_index_4_share, output_sum_secondmodule_equation_num_5_index_5_share, output_sum_secondmodule_equation_num_5_index_6_share, output_sum_secondmodule_equation_num_5_index_7_share, output_sum_secondmodule_equation_num_5_index_8_share, output_sum_secondmodule_equation_num_5_index_9_share, output_sum_secondmodule_equation_num_5_index_10_share, output_sum_secondmodule_equation_num_5_index_11_share, output_sum_secondmodule_equation_num_5_index_12_share, output_sum_secondmodule_equation_num_5_index_13_share, output_sum_secondmodule_equation_num_5_index_14_share;
output output_sum_secondmodule_equation_num_6_index_0_share, output_sum_secondmodule_equation_num_6_index_1_share, output_sum_secondmodule_equation_num_6_index_2_share, output_sum_secondmodule_equation_num_6_index_3_share, output_sum_secondmodule_equation_num_6_index_4_share, output_sum_secondmodule_equation_num_6_index_5_share, output_sum_secondmodule_equation_num_6_index_6_share, output_sum_secondmodule_equation_num_6_index_7_share, output_sum_secondmodule_equation_num_6_index_8_share, output_sum_secondmodule_equation_num_6_index_9_share, output_sum_secondmodule_equation_num_6_index_10_share, output_sum_secondmodule_equation_num_6_index_11_share, output_sum_secondmodule_equation_num_6_index_12_share, output_sum_secondmodule_equation_num_6_index_13_share, output_sum_secondmodule_equation_num_6_index_14_share;
output output_sum_secondmodule_equation_num_7_index_0_share, output_sum_secondmodule_equation_num_7_index_1_share, output_sum_secondmodule_equation_num_7_index_2_share, output_sum_secondmodule_equation_num_7_index_3_share, output_sum_secondmodule_equation_num_7_index_4_share, output_sum_secondmodule_equation_num_7_index_5_share, output_sum_secondmodule_equation_num_7_index_6_share, output_sum_secondmodule_equation_num_7_index_7_share, output_sum_secondmodule_equation_num_7_index_8_share, output_sum_secondmodule_equation_num_7_index_9_share, output_sum_secondmodule_equation_num_7_index_10_share, output_sum_secondmodule_equation_num_7_index_11_share, output_sum_secondmodule_equation_num_7_index_12_share, output_sum_secondmodule_equation_num_7_index_13_share, output_sum_secondmodule_equation_num_7_index_14_share;




assign output_sum_secondmodule_equation_num_0_index_0_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_1_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_2_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_3_share =  ( ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_4_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_5_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_6_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_7_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_8_share =  ( ( output_x4_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_9_share =  ( ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_10_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_11_share =  ( ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_12_share =  ( ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_13_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_0_index_14_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x6x7_share ) ) ;




assign output_sum_secondmodule_equation_num_1_index_0_share =  ( ( output_x4_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_1_share =  ( ( output_x4_share ) ^ ( output_x7_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_2_share =  ( ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_3_share =  ( ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_4_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_5_share =  ( ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_6_share =  ( ( output_x4_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_7_share =  ( ( output_x4_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_8_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_9_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_10_share =  ( ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_11_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_12_share =  ( ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_13_share =  ( ( output_x5_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_1_index_14_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;




assign output_sum_secondmodule_equation_num_2_index_0_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_1_share =  ( ( output_x4_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_2_share =  ( ( output_x4x5_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_3_share =  ( ( output_x4_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_4_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_5_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_6_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_7_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_8_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_9_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_10_share =  ( ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_11_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_12_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_13_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_2_index_14_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;




assign output_sum_secondmodule_equation_num_3_index_0_share =  ( ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_1_share =  ( ( output_x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_2_share =  ( ( output_x4x5_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_3_share =  ( ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_4_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_5_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_6_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_7_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_8_share =  ( ( output_x4_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_9_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_10_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_11_share =  ( ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_12_share =  ( ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_13_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_3_index_14_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ) ;




assign output_sum_secondmodule_equation_num_4_index_0_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_1_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_2_share =  ( ( output_x5_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_3_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_4_share =  ( ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_5_share =  ( ( output_x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_6_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_7_share =  ( ( output_x4_share ) ^ ( output_x4x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_8_share =  ( ( output_x5_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_9_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_10_share =  ( ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_11_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_12_share =  ( ( output_x4_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_13_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_4_index_14_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;


assign output_sum_secondmodule_equation_num_5_index_0_share =  ( ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_1_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_2_share =  ( ( output_x4_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_3_share =  ( ( output_x4_share ) ^ ( output_x4x5_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_4_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_5_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_6_share =  ( ( output_x5_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_7_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_8_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_9_share =  ( ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_10_share =  ( ( output_x5_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_11_share =  ( ( output_x4_share ) ^ ( output_x7_share ) ^ ( output_x5x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_12_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_13_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_5_index_14_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x5x6x7_share ) ) ;



assign output_sum_secondmodule_equation_num_6_index_0_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_1_share =  ( ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_2_share =  ( ( output_x4x6_share ) ^ ( output_x4x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_3_share =  ( ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_4_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_5_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_6_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_7_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_8_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_9_share =  ( ( output_x4_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_10_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_11_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_12_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x5x6_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_13_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x5x7_share ) ) ;
assign output_sum_secondmodule_equation_num_6_index_14_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ) ;



assign output_sum_secondmodule_equation_num_7_index_0_share =  ( ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x5x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_1_share =  ( ( output_x7_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_2_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x4x6_share ) ^ ( output_x5x6_share ) ^ ( output_x6x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_3_share =  ( ( output_x5_share ) ^ ( output_x4x5_share ) ^ ( output_x5x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_4_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_5_share =  ( ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_6_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x5x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_7_share =  ( ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_8_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x4x7_share ) ^ ( output_x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_9_share =  ( ( output_x5_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_10_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x4x6_share ) ^ ( output_x5x7_share ) ^ ( output_x6x7_share ) ^ ( output_x4x5x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_11_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x4x5_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_12_share =  ( ( output_x5_share ) ^ ( output_x6_share ) ^ ( output_x7_share ) ^ ( output_x4x5_share ) ^ ( output_x4x6_share ) ^ ( output_x4x7_share ) ^ ( output_x4x5x6_share ) ^ ( output_x4x5x7_share ) ^ ( output_x4x6x7_share ) ^ ( output_x5x6x7_share ) ^ ( output_x4x5x6x7_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_13_share =  ( ( output_x4_share ) ^ ( output_x5_share ) ^ ( output_x7_share ) ^ ( output_x5x6_share ) ) ;
assign output_sum_secondmodule_equation_num_7_index_14_share =  ( ( output_x4_share ) ^ ( output_x6_share ) ^ ( output_x6x7_share ) ) ;

endmodule