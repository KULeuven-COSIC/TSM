`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 22:00:00 02/22/2025
// Design Name: Second-Order Masked AES S-Box
// Module Name: AES_sbox_secondorder_tworegstages_final
// Project Name: PINI Second-Order Two-Cycle AES S-Box
// Target Device: FPGA
// Tool Version: Vivado 2020.2
// Description: Implements a second-order masked AES S-Box using HO-TSM with two register stages.
// Dependencies: None
//
// Revision:
// Revision 0.02 - Optimized combinatorial logic for two-cycle computation
////////////////////////////////////////////////////////////////////////////////

module AES_sbox_secondorder_tworegstages_final ( 
    clk, 
    rand_bit_cycle1, rand_bit_cycle2,
	sbox_input_share1, sbox_input_share2, sbox_input_share3,
    output_share1, output_share2, output_share3
);


input clk;

input [278:1] rand_bit_cycle1;
input [508:1] rand_bit_cycle2;

input [7:0] sbox_input_share1, sbox_input_share2, sbox_input_share3;
output [7:0] output_share1, output_share2, output_share3;

wire [8:1] rand_composable_bit_a;
wire [8:1] rand_composable_bit_b;
wire [8:1] rand_composable_bit_c;

assign rand_composable_bit_a = rand_bit_cycle1[8:1] ;
assign rand_composable_bit_b = rand_bit_cycle1[16:9] ;
assign rand_composable_bit_c = rand_bit_cycle1[24:17] ;

wire x0_input_share1 = sbox_input_share1[0] ^ rand_composable_bit_a[1] ^ rand_composable_bit_c[1] ;
wire x1_input_share1 = sbox_input_share1[1] ^ rand_composable_bit_a[2] ^ rand_composable_bit_c[2] ;
wire x2_input_share1 = sbox_input_share1[2] ^ rand_composable_bit_a[3] ^ rand_composable_bit_c[3] ;
wire x3_input_share1 = sbox_input_share1[3] ^ rand_composable_bit_a[4] ^ rand_composable_bit_c[4] ;
wire x4_input_share1 = sbox_input_share1[4] ^ rand_composable_bit_a[5] ^ rand_composable_bit_c[5] ;
wire x5_input_share1 = sbox_input_share1[5] ^ rand_composable_bit_a[6] ^ rand_composable_bit_c[6] ;
wire x6_input_share1 = sbox_input_share1[6] ^ rand_composable_bit_a[7] ^ rand_composable_bit_c[7] ;
wire x7_input_share1 = sbox_input_share1[7] ^ rand_composable_bit_a[8] ^ rand_composable_bit_c[8] ;

wire x0_input_share2 = sbox_input_share2[0] ^ rand_composable_bit_b[1] ^ rand_composable_bit_c[1] ;
wire x1_input_share2 = sbox_input_share2[1] ^ rand_composable_bit_b[2] ^ rand_composable_bit_c[2] ;
wire x2_input_share2 = sbox_input_share2[2] ^ rand_composable_bit_b[3] ^ rand_composable_bit_c[3] ;
wire x3_input_share2 = sbox_input_share2[3] ^ rand_composable_bit_b[4] ^ rand_composable_bit_c[4] ;
wire x4_input_share2 = sbox_input_share2[4] ^ rand_composable_bit_b[5] ^ rand_composable_bit_c[5] ;
wire x5_input_share2 = sbox_input_share2[5] ^ rand_composable_bit_b[6] ^ rand_composable_bit_c[6] ;
wire x6_input_share2 = sbox_input_share2[6] ^ rand_composable_bit_b[7] ^ rand_composable_bit_c[7] ;
wire x7_input_share2 = sbox_input_share2[7] ^ rand_composable_bit_b[8] ^ rand_composable_bit_c[8] ;

wire x0_input_share3 = sbox_input_share3[0] ^ rand_composable_bit_a[1]  ^ rand_composable_bit_b[1] ;
wire x1_input_share3 = sbox_input_share3[1] ^ rand_composable_bit_a[2]  ^ rand_composable_bit_b[2] ;
wire x2_input_share3 = sbox_input_share3[2] ^ rand_composable_bit_a[3]  ^ rand_composable_bit_b[3] ;
wire x3_input_share3 = sbox_input_share3[3] ^ rand_composable_bit_a[4]  ^ rand_composable_bit_b[4] ;
wire x4_input_share3 = sbox_input_share3[4] ^ rand_composable_bit_a[5]  ^ rand_composable_bit_b[5] ;
wire x5_input_share3 = sbox_input_share3[5] ^ rand_composable_bit_a[6]  ^ rand_composable_bit_b[6] ;
wire x6_input_share3 = sbox_input_share3[6] ^ rand_composable_bit_a[7]  ^ rand_composable_bit_b[7] ;
wire x7_input_share3 = sbox_input_share3[7] ^ rand_composable_bit_a[8]  ^ rand_composable_bit_b[8] ;



// Cycle 1 Logic

allcrossproducts_oneshare_eightinputs first_cycle(
x0_input_share1 ,x1_input_share1 ,x2_input_share1 ,x3_input_share1 ,x4_input_share1 ,x5_input_share1 ,x6_input_share1 ,x7_input_share1 ,
x0_subscript0_sharex             , x1_subscript0_sharex             , x2_subscript0_sharex             , x3_subscript0_sharex             , x4_subscript0_sharex             , x5_subscript0_sharex             , x6_subscript0_sharex             , x7_subscript0_sharex             , x0x1_subscript0_sharex           , x0x4_subscript0_sharex           , x0x5_subscript0_sharex           , x0x6_subscript0_sharex           , x1x2_subscript0_sharex           , x1x3_subscript0_sharex           , x1x4_subscript0_sharex           , x1x6_subscript0_sharex           , x2x3_subscript0_sharex           , x2x4_subscript0_sharex           , x2x6_subscript0_sharex           , x2x7_subscript0_sharex           , x4x6_subscript0_sharex           , x5x6_subscript0_sharex           , x5x7_subscript0_sharex           , x6x7_subscript0_sharex           , x0x2_subscript0_sharex           , x0x3_subscript0_sharex           , x0x7_subscript0_sharex           , x1x7_subscript0_sharex           , x3x7_subscript0_sharex           , x4x5_subscript0_sharex           , x3x4_subscript0_sharex           , x4x7_subscript0_sharex           , x3x6_subscript0_sharex           , x1x5_subscript0_sharex           , x2x5_subscript0_sharex           , x3x5_subscript0_sharex           , x0x1x4_subscript0_sharex         , x0x1x6_subscript0_sharex         , x0x1x7_subscript0_sharex         , x0x2x4_subscript0_sharex         , x0x2x5_subscript0_sharex         , x0x2x6_subscript0_sharex         , x0x2x7_subscript0_sharex         , x0x3x4_subscript0_sharex         , x0x3x5_subscript0_sharex         , x0x3x6_subscript0_sharex         , x0x4x6_subscript0_sharex         , x0x4x7_subscript0_sharex         , x1x2x3_subscript0_sharex         , x1x2x4_subscript0_sharex         , x1x2x6_subscript0_sharex         , x1x3x4_subscript0_sharex         , x1x3x7_subscript0_sharex         , x1x4x6_subscript0_sharex         , x1x5x6_subscript0_sharex         , x2x3x5_subscript0_sharex         , x2x3x7_subscript0_sharex         , x2x4x7_subscript0_sharex         , x2x5x6_subscript0_sharex         , x2x5x7_subscript0_sharex         , x2x6x7_subscript0_sharex         , x3x4x7_subscript0_sharex         , x3x5x7_subscript0_sharex         , x3x6x7_subscript0_sharex         , x4x5x6_subscript0_sharex         , x5x6x7_subscript0_sharex         , x0x1x3_subscript0_sharex         , x0x2x3_subscript0_sharex         , x0x4x5_subscript0_sharex         , x0x5x7_subscript0_sharex         , x0x6x7_subscript0_sharex         , x1x3x5_subscript0_sharex         , x1x3x6_subscript0_sharex         , x1x4x7_subscript0_sharex         , x2x3x4_subscript0_sharex         , x2x3x6_subscript0_sharex         , x3x4x6_subscript0_sharex         , x3x5x6_subscript0_sharex         , x0x1x5_subscript0_sharex         , x0x3x7_subscript0_sharex         , x1x2x5_subscript0_sharex         , x1x2x7_subscript0_sharex         , x1x4x5_subscript0_sharex         , x1x5x7_subscript0_sharex         , x2x4x5_subscript0_sharex         , x3x4x5_subscript0_sharex         , x4x6x7_subscript0_sharex         , x1x6x7_subscript0_sharex         , x4x5x7_subscript0_sharex         , x0x1x2_subscript0_sharex         , x0x5x6_subscript0_sharex         , x2x4x6_subscript0_sharex         , x0x1x2x3_subscript0_sharex       , x0x1x2x5_subscript0_sharex       , x0x1x2x6_subscript0_sharex       , x0x1x2x7_subscript0_sharex       , x0x1x4x5_subscript0_sharex       , x0x1x4x7_subscript0_sharex       , x0x2x3x5_subscript0_sharex       , x0x2x3x7_subscript0_sharex       , x0x2x4x5_subscript0_sharex       , x0x2x4x7_subscript0_sharex       , x0x2x5x6_subscript0_sharex       , x0x2x5x7_subscript0_sharex       , x0x3x4x6_subscript0_sharex       , x0x3x5x6_subscript0_sharex       , x0x4x5x6_subscript0_sharex       , x0x4x5x7_subscript0_sharex       , x0x4x6x7_subscript0_sharex       , x1x2x3x5_subscript0_sharex       , x1x2x3x6_subscript0_sharex       , x1x2x3x7_subscript0_sharex       , x1x2x4x6_subscript0_sharex       , x1x2x4x7_subscript0_sharex       , x1x2x6x7_subscript0_sharex       , x1x3x4x6_subscript0_sharex       , x1x3x6x7_subscript0_sharex       , x1x4x5x6_subscript0_sharex       , x1x4x5x7_subscript0_sharex       , x1x5x6x7_subscript0_sharex       , x2x3x5x7_subscript0_sharex       , x2x3x6x7_subscript0_sharex       , x2x4x5x6_subscript0_sharex       , x2x4x5x7_subscript0_sharex       , x3x5x6x7_subscript0_sharex       , x0x1x3x4_subscript0_sharex       , x0x1x3x6_subscript0_sharex       , x0x1x5x6_subscript0_sharex       , x0x2x3x6_subscript0_sharex       , x0x3x4x5_subscript0_sharex       , x1x2x5x6_subscript0_sharex       , x1x2x5x7_subscript0_sharex       , x1x3x4x5_subscript0_sharex       , x1x3x4x7_subscript0_sharex       , x1x3x5x6_subscript0_sharex       , x1x3x5x7_subscript0_sharex       , x1x4x6x7_subscript0_sharex       , x2x3x4x5_subscript0_sharex       , x2x3x4x7_subscript0_sharex       , x2x4x6x7_subscript0_sharex       , x3x4x5x6_subscript0_sharex       , x3x4x5x7_subscript0_sharex       , x3x4x6x7_subscript0_sharex       , x0x1x3x5_subscript0_sharex       , x0x1x4x6_subscript0_sharex       , x0x2x3x4_subscript0_sharex       , x0x2x4x6_subscript0_sharex       , x0x3x4x7_subscript0_sharex       , x0x3x5x7_subscript0_sharex       , x1x2x3x4_subscript0_sharex       , x2x3x4x6_subscript0_sharex       , x2x3x5x6_subscript0_sharex       , x2x5x6x7_subscript0_sharex       , x4x5x6x7_subscript0_sharex       , x0x1x2x4_subscript0_sharex       , x0x1x6x7_subscript0_sharex       , x0x2x6x7_subscript0_sharex       , x0x3x6x7_subscript0_sharex       , x0x5x6x7_subscript0_sharex       , x1x2x4x5_subscript0_sharex       , x0x1x3x7_subscript0_sharex       , x0x1x5x7_subscript0_sharex       , x0x1x2x3x4_subscript0_sharex     , x0x1x2x3x6_subscript0_sharex     , x0x1x2x3x7_subscript0_sharex     , x0x1x2x4x5_subscript0_sharex     , x0x1x2x4x7_subscript0_sharex     , x0x1x2x5x7_subscript0_sharex     , x0x1x2x6x7_subscript0_sharex     , x0x1x3x4x6_subscript0_sharex     , x0x1x3x5x6_subscript0_sharex     , x0x1x3x5x7_subscript0_sharex     , x0x1x3x6x7_subscript0_sharex     , x0x1x4x5x6_subscript0_sharex     , x0x1x5x6x7_subscript0_sharex     , x0x2x3x4x5_subscript0_sharex     , x0x2x3x4x6_subscript0_sharex     , x0x2x4x5x7_subscript0_sharex     , x0x2x4x6x7_subscript0_sharex     , x0x3x4x5x6_subscript0_sharex     , x0x3x4x5x7_subscript0_sharex     , x0x3x4x6x7_subscript0_sharex     , x0x3x5x6x7_subscript0_sharex     , x1x2x3x5x6_subscript0_sharex     , x1x2x3x5x7_subscript0_sharex     , x1x2x4x5x6_subscript0_sharex     , x1x2x4x6x7_subscript0_sharex     , x1x2x5x6x7_subscript0_sharex     , x1x3x4x5x7_subscript0_sharex     , x2x3x4x5x6_subscript0_sharex     , x2x3x4x5x7_subscript0_sharex     , x2x4x5x6x7_subscript0_sharex     , x0x1x2x4x6_subscript0_sharex     , x0x1x3x4x7_subscript0_sharex     , x0x2x3x4x7_subscript0_sharex     , x0x2x3x5x7_subscript0_sharex     , x0x2x3x6x7_subscript0_sharex     , x0x2x4x5x6_subscript0_sharex     , x0x2x5x6x7_subscript0_sharex     , x0x4x5x6x7_subscript0_sharex     , x1x2x3x4x6_subscript0_sharex     , x1x3x4x5x6_subscript0_sharex     , x2x3x4x6x7_subscript0_sharex     , x0x1x2x3x5_subscript0_sharex     , x0x1x4x6x7_subscript0_sharex     , x1x2x3x4x5_subscript0_sharex     , x1x2x3x6x7_subscript0_sharex     , x1x2x4x5x7_subscript0_sharex     , x1x3x4x6x7_subscript0_sharex     , x1x3x5x6x7_subscript0_sharex     , x1x4x5x6x7_subscript0_sharex     , x2x3x5x6x7_subscript0_sharex     , x3x4x5x6x7_subscript0_sharex     , x0x1x2x5x6_subscript0_sharex     , x0x1x3x4x5_subscript0_sharex     , x0x1x4x5x7_subscript0_sharex     , x0x2x3x5x6_subscript0_sharex     , x1x2x3x4x7_subscript0_sharex     , x0x1x2x3x4x6_subscript0_sharex   , x0x1x2x3x4x7_subscript0_sharex   , x0x1x2x3x5x7_subscript0_sharex   , x0x1x2x3x6x7_subscript0_sharex   , x0x1x2x4x5x7_subscript0_sharex   , x0x1x2x5x6x7_subscript0_sharex   , x0x1x3x4x6x7_subscript0_sharex   , x0x1x4x5x6x7_subscript0_sharex   , x0x2x3x4x5x6_subscript0_sharex   , x0x2x3x4x5x7_subscript0_sharex   , x0x2x3x5x6x7_subscript0_sharex   , x1x2x3x4x6x7_subscript0_sharex   , x1x2x4x5x6x7_subscript0_sharex   , x1x3x4x5x6x7_subscript0_sharex   , x2x3x4x5x6x7_subscript0_sharex   , x0x1x2x3x5x6_subscript0_sharex   , x0x1x2x4x6x7_subscript0_sharex   , x0x1x3x4x5x6_subscript0_sharex   , x0x2x3x4x6x7_subscript0_sharex   , x1x2x3x4x5x6_subscript0_sharex   , x1x2x3x5x6x7_subscript0_sharex   , x0x1x2x3x4x5_subscript0_sharex   , x0x1x2x4x5x6_subscript0_sharex   , x0x1x3x4x5x7_subscript0_sharex   , x0x1x3x5x6x7_subscript0_sharex   , x0x2x4x5x6x7_subscript0_sharex   , x1x2x3x4x5x7_subscript0_sharex   , x0x3x4x5x6x7_subscript0_sharex   , x0x1x2x3x4x6x7_subscript0_sharex , x0x1x2x4x5x6x7_subscript0_sharex , x0x2x3x4x5x6x7_subscript0_sharex , x0x1x2x3x5x6x7_subscript0_sharex , x0x1x3x4x5x6x7_subscript0_sharex , x1x2x3x4x5x6x7_subscript0_sharex , x0x1x2x3x4x5x6_subscript0_sharex , x0x1x2x3x4x5x7_subscript0_sharex
);

wire [254:1] rand_first_cycle ;
assign rand_first_cycle = rand_bit_cycle1[278:25];

xor_AES_twofiftyfour first_cycle_xor(
x0_subscript0_sharex             , x1_subscript0_sharex             , x2_subscript0_sharex             , x3_subscript0_sharex             , x4_subscript0_sharex             , x5_subscript0_sharex             , x6_subscript0_sharex             , x7_subscript0_sharex             , x0x1_subscript0_sharex           , x0x4_subscript0_sharex           , x0x5_subscript0_sharex           , x0x6_subscript0_sharex           , x1x2_subscript0_sharex           , x1x3_subscript0_sharex           , x1x4_subscript0_sharex           , x1x6_subscript0_sharex           , x2x3_subscript0_sharex           , x2x4_subscript0_sharex           , x2x6_subscript0_sharex           , x2x7_subscript0_sharex           , x4x6_subscript0_sharex           , x5x6_subscript0_sharex           , x5x7_subscript0_sharex           , x6x7_subscript0_sharex           , x0x2_subscript0_sharex           , x0x3_subscript0_sharex           , x0x7_subscript0_sharex           , x1x7_subscript0_sharex           , x3x7_subscript0_sharex           , x4x5_subscript0_sharex           , x3x4_subscript0_sharex           , x4x7_subscript0_sharex           , x3x6_subscript0_sharex           , x1x5_subscript0_sharex           , x2x5_subscript0_sharex           , x3x5_subscript0_sharex           , x0x1x4_subscript0_sharex         , x0x1x6_subscript0_sharex         , x0x1x7_subscript0_sharex         , x0x2x4_subscript0_sharex         , x0x2x5_subscript0_sharex         , x0x2x6_subscript0_sharex         , x0x2x7_subscript0_sharex         , x0x3x4_subscript0_sharex         , x0x3x5_subscript0_sharex         , x0x3x6_subscript0_sharex         , x0x4x6_subscript0_sharex         , x0x4x7_subscript0_sharex         , x1x2x3_subscript0_sharex         , x1x2x4_subscript0_sharex         , x1x2x6_subscript0_sharex         , x1x3x4_subscript0_sharex         , x1x3x7_subscript0_sharex         , x1x4x6_subscript0_sharex         , x1x5x6_subscript0_sharex         , x2x3x5_subscript0_sharex         , x2x3x7_subscript0_sharex         , x2x4x7_subscript0_sharex         , x2x5x6_subscript0_sharex         , x2x5x7_subscript0_sharex         , x2x6x7_subscript0_sharex         , x3x4x7_subscript0_sharex         , x3x5x7_subscript0_sharex         , x3x6x7_subscript0_sharex         , x4x5x6_subscript0_sharex         , x5x6x7_subscript0_sharex         , x0x1x3_subscript0_sharex         , x0x2x3_subscript0_sharex         , x0x4x5_subscript0_sharex         , x0x5x7_subscript0_sharex         , x0x6x7_subscript0_sharex         , x1x3x5_subscript0_sharex         , x1x3x6_subscript0_sharex         , x1x4x7_subscript0_sharex         , x2x3x4_subscript0_sharex         , x2x3x6_subscript0_sharex         , x3x4x6_subscript0_sharex         , x3x5x6_subscript0_sharex         , x0x1x5_subscript0_sharex         , x0x3x7_subscript0_sharex         , x1x2x5_subscript0_sharex         , x1x2x7_subscript0_sharex         , x1x4x5_subscript0_sharex         , x1x5x7_subscript0_sharex         , x2x4x5_subscript0_sharex         , x3x4x5_subscript0_sharex         , x4x6x7_subscript0_sharex         , x1x6x7_subscript0_sharex         , x4x5x7_subscript0_sharex         , x0x1x2_subscript0_sharex         , x0x5x6_subscript0_sharex         , x2x4x6_subscript0_sharex         , x0x1x2x3_subscript0_sharex       , x0x1x2x5_subscript0_sharex       , x0x1x2x6_subscript0_sharex       , x0x1x2x7_subscript0_sharex       , x0x1x4x5_subscript0_sharex       , x0x1x4x7_subscript0_sharex       , x0x2x3x5_subscript0_sharex       , x0x2x3x7_subscript0_sharex       , x0x2x4x5_subscript0_sharex       , x0x2x4x7_subscript0_sharex       , x0x2x5x6_subscript0_sharex       , x0x2x5x7_subscript0_sharex       , x0x3x4x6_subscript0_sharex       , x0x3x5x6_subscript0_sharex       , x0x4x5x6_subscript0_sharex       , x0x4x5x7_subscript0_sharex       , x0x4x6x7_subscript0_sharex       , x1x2x3x5_subscript0_sharex       , x1x2x3x6_subscript0_sharex       , x1x2x3x7_subscript0_sharex       , x1x2x4x6_subscript0_sharex       , x1x2x4x7_subscript0_sharex       , x1x2x6x7_subscript0_sharex       , x1x3x4x6_subscript0_sharex       , x1x3x6x7_subscript0_sharex       , x1x4x5x6_subscript0_sharex       , x1x4x5x7_subscript0_sharex       , x1x5x6x7_subscript0_sharex       , x2x3x5x7_subscript0_sharex       , x2x3x6x7_subscript0_sharex       , x2x4x5x6_subscript0_sharex       , x2x4x5x7_subscript0_sharex       , x3x5x6x7_subscript0_sharex       , x0x1x3x4_subscript0_sharex       , x0x1x3x6_subscript0_sharex       , x0x1x5x6_subscript0_sharex       , x0x2x3x6_subscript0_sharex       , x0x3x4x5_subscript0_sharex       , x1x2x5x6_subscript0_sharex       , x1x2x5x7_subscript0_sharex       , x1x3x4x5_subscript0_sharex       , x1x3x4x7_subscript0_sharex       , x1x3x5x6_subscript0_sharex       , x1x3x5x7_subscript0_sharex       , x1x4x6x7_subscript0_sharex       , x2x3x4x5_subscript0_sharex       , x2x3x4x7_subscript0_sharex       , x2x4x6x7_subscript0_sharex       , x3x4x5x6_subscript0_sharex       , x3x4x5x7_subscript0_sharex       , x3x4x6x7_subscript0_sharex       , x0x1x3x5_subscript0_sharex       , x0x1x4x6_subscript0_sharex       , x0x2x3x4_subscript0_sharex       , x0x2x4x6_subscript0_sharex       , x0x3x4x7_subscript0_sharex       , x0x3x5x7_subscript0_sharex       , x1x2x3x4_subscript0_sharex       , x2x3x4x6_subscript0_sharex       , x2x3x5x6_subscript0_sharex       , x2x5x6x7_subscript0_sharex       , x4x5x6x7_subscript0_sharex       , x0x1x2x4_subscript0_sharex       , x0x1x6x7_subscript0_sharex       , x0x2x6x7_subscript0_sharex       , x0x3x6x7_subscript0_sharex       , x0x5x6x7_subscript0_sharex       , x1x2x4x5_subscript0_sharex       , x0x1x3x7_subscript0_sharex       , x0x1x5x7_subscript0_sharex       , x0x1x2x3x4_subscript0_sharex     , x0x1x2x3x6_subscript0_sharex     , x0x1x2x3x7_subscript0_sharex     , x0x1x2x4x5_subscript0_sharex     , x0x1x2x4x7_subscript0_sharex     , x0x1x2x5x7_subscript0_sharex     , x0x1x2x6x7_subscript0_sharex     , x0x1x3x4x6_subscript0_sharex     , x0x1x3x5x6_subscript0_sharex     , x0x1x3x5x7_subscript0_sharex     , x0x1x3x6x7_subscript0_sharex     , x0x1x4x5x6_subscript0_sharex     , x0x1x5x6x7_subscript0_sharex     , x0x2x3x4x5_subscript0_sharex     , x0x2x3x4x6_subscript0_sharex     , x0x2x4x5x7_subscript0_sharex     , x0x2x4x6x7_subscript0_sharex     , x0x3x4x5x6_subscript0_sharex     , x0x3x4x5x7_subscript0_sharex     , x0x3x4x6x7_subscript0_sharex     , x0x3x5x6x7_subscript0_sharex     , x1x2x3x5x6_subscript0_sharex     , x1x2x3x5x7_subscript0_sharex     , x1x2x4x5x6_subscript0_sharex     , x1x2x4x6x7_subscript0_sharex     , x1x2x5x6x7_subscript0_sharex     , x1x3x4x5x7_subscript0_sharex     , x2x3x4x5x6_subscript0_sharex     , x2x3x4x5x7_subscript0_sharex     , x2x4x5x6x7_subscript0_sharex     , x0x1x2x4x6_subscript0_sharex     , x0x1x3x4x7_subscript0_sharex     , x0x2x3x4x7_subscript0_sharex     , x0x2x3x5x7_subscript0_sharex     , x0x2x3x6x7_subscript0_sharex     , x0x2x4x5x6_subscript0_sharex     , x0x2x5x6x7_subscript0_sharex     , x0x4x5x6x7_subscript0_sharex     , x1x2x3x4x6_subscript0_sharex     , x1x3x4x5x6_subscript0_sharex     , x2x3x4x6x7_subscript0_sharex     , x0x1x2x3x5_subscript0_sharex     , x0x1x4x6x7_subscript0_sharex     , x1x2x3x4x5_subscript0_sharex     , x1x2x3x6x7_subscript0_sharex     , x1x2x4x5x7_subscript0_sharex     , x1x3x4x6x7_subscript0_sharex     , x1x3x5x6x7_subscript0_sharex     , x1x4x5x6x7_subscript0_sharex     , x2x3x5x6x7_subscript0_sharex     , x3x4x5x6x7_subscript0_sharex     , x0x1x2x5x6_subscript0_sharex     , x0x1x3x4x5_subscript0_sharex     , x0x1x4x5x7_subscript0_sharex     , x0x2x3x5x6_subscript0_sharex     , x1x2x3x4x7_subscript0_sharex     , x0x1x2x3x4x6_subscript0_sharex   , x0x1x2x3x4x7_subscript0_sharex   , x0x1x2x3x5x7_subscript0_sharex   , x0x1x2x3x6x7_subscript0_sharex   , x0x1x2x4x5x7_subscript0_sharex   , x0x1x2x5x6x7_subscript0_sharex   , x0x1x3x4x6x7_subscript0_sharex   , x0x1x4x5x6x7_subscript0_sharex   , x0x2x3x4x5x6_subscript0_sharex   , x0x2x3x4x5x7_subscript0_sharex   , x0x2x3x5x6x7_subscript0_sharex   , x1x2x3x4x6x7_subscript0_sharex   , x1x2x4x5x6x7_subscript0_sharex   , x1x3x4x5x6x7_subscript0_sharex   , x2x3x4x5x6x7_subscript0_sharex   , x0x1x2x3x5x6_subscript0_sharex   , x0x1x2x4x6x7_subscript0_sharex   , x0x1x3x4x5x6_subscript0_sharex   , x0x2x3x4x6x7_subscript0_sharex   , x1x2x3x4x5x6_subscript0_sharex   , x1x2x3x5x6x7_subscript0_sharex   , x0x1x2x3x4x5_subscript0_sharex   , x0x1x2x4x5x6_subscript0_sharex   , x0x1x3x4x5x7_subscript0_sharex   , x0x1x3x5x6x7_subscript0_sharex   , x0x2x4x5x6x7_subscript0_sharex   , x1x2x3x4x5x7_subscript0_sharex   , x0x3x4x5x6x7_subscript0_sharex   , x0x1x2x3x4x6x7_subscript0_sharex , x0x1x2x4x5x6x7_subscript0_sharex , x0x2x3x4x5x6x7_subscript0_sharex , x0x1x2x3x5x6x7_subscript0_sharex , x0x1x3x4x5x6x7_subscript0_sharex , x1x2x3x4x5x6x7_subscript0_sharex , x0x1x2x3x4x5x6_subscript0_sharex , x0x1x2x3x4x5x7_subscript0_sharex ,
rand_first_cycle[1] ,rand_first_cycle[2] ,rand_first_cycle[3] ,rand_first_cycle[4] ,rand_first_cycle[5] ,rand_first_cycle[6] ,rand_first_cycle[7] ,rand_first_cycle[8] ,rand_first_cycle[9] ,rand_first_cycle[10] ,rand_first_cycle[11] ,rand_first_cycle[12] ,rand_first_cycle[13] ,rand_first_cycle[14] ,rand_first_cycle[15] ,rand_first_cycle[16] ,rand_first_cycle[17] ,rand_first_cycle[18] ,rand_first_cycle[19] ,rand_first_cycle[20] ,rand_first_cycle[21] ,rand_first_cycle[22] ,rand_first_cycle[23] ,rand_first_cycle[24] ,rand_first_cycle[25] ,rand_first_cycle[26] ,rand_first_cycle[27] ,rand_first_cycle[28] ,rand_first_cycle[29] ,rand_first_cycle[30] ,rand_first_cycle[31] ,rand_first_cycle[32] ,rand_first_cycle[33] ,rand_first_cycle[34] ,rand_first_cycle[35] ,rand_first_cycle[36] ,rand_first_cycle[37] ,rand_first_cycle[38] ,rand_first_cycle[39] ,rand_first_cycle[40] ,rand_first_cycle[41] ,rand_first_cycle[42] ,rand_first_cycle[43] ,rand_first_cycle[44] ,rand_first_cycle[45] ,rand_first_cycle[46] ,rand_first_cycle[47] ,rand_first_cycle[48] ,rand_first_cycle[49] ,rand_first_cycle[50] ,rand_first_cycle[51] ,rand_first_cycle[52] ,rand_first_cycle[53] ,rand_first_cycle[54] ,rand_first_cycle[55] ,rand_first_cycle[56] ,rand_first_cycle[57] ,rand_first_cycle[58] ,rand_first_cycle[59] ,rand_first_cycle[60] ,rand_first_cycle[61] ,rand_first_cycle[62] ,rand_first_cycle[63] ,rand_first_cycle[64] ,rand_first_cycle[65] ,rand_first_cycle[66] ,rand_first_cycle[67] ,rand_first_cycle[68] ,rand_first_cycle[69] ,rand_first_cycle[70] ,rand_first_cycle[71] ,rand_first_cycle[72] ,rand_first_cycle[73] ,rand_first_cycle[74] ,rand_first_cycle[75] ,rand_first_cycle[76] ,rand_first_cycle[77] ,rand_first_cycle[78] ,rand_first_cycle[79] ,rand_first_cycle[80] ,rand_first_cycle[81] ,rand_first_cycle[82] ,rand_first_cycle[83] ,rand_first_cycle[84] ,rand_first_cycle[85] ,rand_first_cycle[86] ,rand_first_cycle[87] ,rand_first_cycle[88] ,rand_first_cycle[89] ,rand_first_cycle[90] ,rand_first_cycle[91] ,rand_first_cycle[92] ,rand_first_cycle[93] ,rand_first_cycle[94] ,rand_first_cycle[95] ,rand_first_cycle[96] ,rand_first_cycle[97] ,rand_first_cycle[98] ,rand_first_cycle[99] ,rand_first_cycle[100] ,rand_first_cycle[101] ,rand_first_cycle[102] ,rand_first_cycle[103] ,rand_first_cycle[104] ,rand_first_cycle[105] ,rand_first_cycle[106] ,rand_first_cycle[107] ,rand_first_cycle[108] ,rand_first_cycle[109] ,rand_first_cycle[110] ,rand_first_cycle[111] ,rand_first_cycle[112] ,rand_first_cycle[113] ,rand_first_cycle[114] ,rand_first_cycle[115] ,rand_first_cycle[116] ,rand_first_cycle[117] ,rand_first_cycle[118] ,rand_first_cycle[119] ,rand_first_cycle[120] ,rand_first_cycle[121] ,rand_first_cycle[122] ,rand_first_cycle[123] ,rand_first_cycle[124] ,rand_first_cycle[125] ,rand_first_cycle[126] ,rand_first_cycle[127] ,rand_first_cycle[128] ,rand_first_cycle[129] ,rand_first_cycle[130] ,rand_first_cycle[131] ,rand_first_cycle[132] ,rand_first_cycle[133] ,rand_first_cycle[134] ,rand_first_cycle[135] ,rand_first_cycle[136] ,rand_first_cycle[137] ,rand_first_cycle[138] ,rand_first_cycle[139] ,rand_first_cycle[140] ,rand_first_cycle[141] ,rand_first_cycle[142] ,rand_first_cycle[143] ,rand_first_cycle[144] ,rand_first_cycle[145] ,rand_first_cycle[146] ,rand_first_cycle[147] ,rand_first_cycle[148] ,rand_first_cycle[149] ,rand_first_cycle[150] ,rand_first_cycle[151] ,rand_first_cycle[152] ,rand_first_cycle[153] ,rand_first_cycle[154] ,rand_first_cycle[155] ,rand_first_cycle[156] ,rand_first_cycle[157] ,rand_first_cycle[158] ,rand_first_cycle[159] ,rand_first_cycle[160] ,rand_first_cycle[161] ,rand_first_cycle[162] ,rand_first_cycle[163] ,rand_first_cycle[164] ,rand_first_cycle[165] ,rand_first_cycle[166] ,rand_first_cycle[167] ,rand_first_cycle[168] ,rand_first_cycle[169] ,rand_first_cycle[170] ,rand_first_cycle[171] ,rand_first_cycle[172] ,rand_first_cycle[173] ,rand_first_cycle[174] ,rand_first_cycle[175] ,rand_first_cycle[176] ,rand_first_cycle[177] ,rand_first_cycle[178] ,rand_first_cycle[179] ,rand_first_cycle[180] ,rand_first_cycle[181] ,rand_first_cycle[182] ,rand_first_cycle[183] ,rand_first_cycle[184] ,rand_first_cycle[185] ,rand_first_cycle[186] ,rand_first_cycle[187] ,rand_first_cycle[188] ,rand_first_cycle[189] ,rand_first_cycle[190] ,rand_first_cycle[191] ,rand_first_cycle[192] ,rand_first_cycle[193] ,rand_first_cycle[194] ,rand_first_cycle[195] ,rand_first_cycle[196] ,rand_first_cycle[197] ,rand_first_cycle[198] ,rand_first_cycle[199] ,rand_first_cycle[200] ,rand_first_cycle[201] ,rand_first_cycle[202] ,rand_first_cycle[203] ,rand_first_cycle[204] ,rand_first_cycle[205] ,rand_first_cycle[206] ,rand_first_cycle[207] ,rand_first_cycle[208] ,rand_first_cycle[209] ,rand_first_cycle[210] ,rand_first_cycle[211] ,rand_first_cycle[212] ,rand_first_cycle[213] ,rand_first_cycle[214] ,rand_first_cycle[215] ,rand_first_cycle[216] ,rand_first_cycle[217] ,rand_first_cycle[218] ,rand_first_cycle[219] ,rand_first_cycle[220] ,rand_first_cycle[221] ,rand_first_cycle[222] ,rand_first_cycle[223] ,rand_first_cycle[224] ,rand_first_cycle[225] ,rand_first_cycle[226] ,rand_first_cycle[227] ,rand_first_cycle[228] ,rand_first_cycle[229] ,rand_first_cycle[230] ,rand_first_cycle[231] ,rand_first_cycle[232] ,rand_first_cycle[233] ,rand_first_cycle[234] ,rand_first_cycle[235] ,rand_first_cycle[236] ,rand_first_cycle[237] ,rand_first_cycle[238] ,rand_first_cycle[239] ,rand_first_cycle[240] ,rand_first_cycle[241] ,rand_first_cycle[242] ,rand_first_cycle[243] ,rand_first_cycle[244] ,rand_first_cycle[245] ,rand_first_cycle[246] ,rand_first_cycle[247] ,rand_first_cycle[248] ,rand_first_cycle[249] ,rand_first_cycle[250] ,rand_first_cycle[251] ,rand_first_cycle[252] ,rand_first_cycle[253] ,rand_first_cycle[254] ,
x0_subscript0_share1             , x1_subscript0_share1             , x2_subscript0_share1             , x3_subscript0_share1             , x4_subscript0_share1             , x5_subscript0_share1             , x6_subscript0_share1             , x7_subscript0_share1             , x0x1_subscript0_share1           , x0x4_subscript0_share1           , x0x5_subscript0_share1           , x0x6_subscript0_share1           , x1x2_subscript0_share1           , x1x3_subscript0_share1           , x1x4_subscript0_share1           , x1x6_subscript0_share1           , x2x3_subscript0_share1           , x2x4_subscript0_share1           , x2x6_subscript0_share1           , x2x7_subscript0_share1           , x4x6_subscript0_share1           , x5x6_subscript0_share1           , x5x7_subscript0_share1           , x6x7_subscript0_share1           , x0x2_subscript0_share1           , x0x3_subscript0_share1           , x0x7_subscript0_share1           , x1x7_subscript0_share1           , x3x7_subscript0_share1           , x4x5_subscript0_share1           , x3x4_subscript0_share1           , x4x7_subscript0_share1           , x3x6_subscript0_share1           , x1x5_subscript0_share1           , x2x5_subscript0_share1           , x3x5_subscript0_share1           , x0x1x4_subscript0_share1         , x0x1x6_subscript0_share1         , x0x1x7_subscript0_share1         , x0x2x4_subscript0_share1         , x0x2x5_subscript0_share1         , x0x2x6_subscript0_share1         , x0x2x7_subscript0_share1         , x0x3x4_subscript0_share1         , x0x3x5_subscript0_share1         , x0x3x6_subscript0_share1         , x0x4x6_subscript0_share1         , x0x4x7_subscript0_share1         , x1x2x3_subscript0_share1         , x1x2x4_subscript0_share1         , x1x2x6_subscript0_share1         , x1x3x4_subscript0_share1         , x1x3x7_subscript0_share1         , x1x4x6_subscript0_share1         , x1x5x6_subscript0_share1         , x2x3x5_subscript0_share1         , x2x3x7_subscript0_share1         , x2x4x7_subscript0_share1         , x2x5x6_subscript0_share1         , x2x5x7_subscript0_share1         , x2x6x7_subscript0_share1         , x3x4x7_subscript0_share1         , x3x5x7_subscript0_share1         , x3x6x7_subscript0_share1         , x4x5x6_subscript0_share1         , x5x6x7_subscript0_share1         , x0x1x3_subscript0_share1         , x0x2x3_subscript0_share1         , x0x4x5_subscript0_share1         , x0x5x7_subscript0_share1         , x0x6x7_subscript0_share1         , x1x3x5_subscript0_share1         , x1x3x6_subscript0_share1         , x1x4x7_subscript0_share1         , x2x3x4_subscript0_share1         , x2x3x6_subscript0_share1         , x3x4x6_subscript0_share1         , x3x5x6_subscript0_share1         , x0x1x5_subscript0_share1         , x0x3x7_subscript0_share1         , x1x2x5_subscript0_share1         , x1x2x7_subscript0_share1         , x1x4x5_subscript0_share1         , x1x5x7_subscript0_share1         , x2x4x5_subscript0_share1         , x3x4x5_subscript0_share1         , x4x6x7_subscript0_share1         , x1x6x7_subscript0_share1         , x4x5x7_subscript0_share1         , x0x1x2_subscript0_share1         , x0x5x6_subscript0_share1         , x2x4x6_subscript0_share1         , x0x1x2x3_subscript0_share1       , x0x1x2x5_subscript0_share1       , x0x1x2x6_subscript0_share1       , x0x1x2x7_subscript0_share1       , x0x1x4x5_subscript0_share1       , x0x1x4x7_subscript0_share1       , x0x2x3x5_subscript0_share1       , x0x2x3x7_subscript0_share1       , x0x2x4x5_subscript0_share1       , x0x2x4x7_subscript0_share1       , x0x2x5x6_subscript0_share1       , x0x2x5x7_subscript0_share1       , x0x3x4x6_subscript0_share1       , x0x3x5x6_subscript0_share1       , x0x4x5x6_subscript0_share1       , x0x4x5x7_subscript0_share1       , x0x4x6x7_subscript0_share1       , x1x2x3x5_subscript0_share1       , x1x2x3x6_subscript0_share1       , x1x2x3x7_subscript0_share1       , x1x2x4x6_subscript0_share1       , x1x2x4x7_subscript0_share1       , x1x2x6x7_subscript0_share1       , x1x3x4x6_subscript0_share1       , x1x3x6x7_subscript0_share1       , x1x4x5x6_subscript0_share1       , x1x4x5x7_subscript0_share1       , x1x5x6x7_subscript0_share1       , x2x3x5x7_subscript0_share1       , x2x3x6x7_subscript0_share1       , x2x4x5x6_subscript0_share1       , x2x4x5x7_subscript0_share1       , x3x5x6x7_subscript0_share1       , x0x1x3x4_subscript0_share1       , x0x1x3x6_subscript0_share1       , x0x1x5x6_subscript0_share1       , x0x2x3x6_subscript0_share1       , x0x3x4x5_subscript0_share1       , x1x2x5x6_subscript0_share1       , x1x2x5x7_subscript0_share1       , x1x3x4x5_subscript0_share1       , x1x3x4x7_subscript0_share1       , x1x3x5x6_subscript0_share1       , x1x3x5x7_subscript0_share1       , x1x4x6x7_subscript0_share1       , x2x3x4x5_subscript0_share1       , x2x3x4x7_subscript0_share1       , x2x4x6x7_subscript0_share1       , x3x4x5x6_subscript0_share1       , x3x4x5x7_subscript0_share1       , x3x4x6x7_subscript0_share1       , x0x1x3x5_subscript0_share1       , x0x1x4x6_subscript0_share1       , x0x2x3x4_subscript0_share1       , x0x2x4x6_subscript0_share1       , x0x3x4x7_subscript0_share1       , x0x3x5x7_subscript0_share1       , x1x2x3x4_subscript0_share1       , x2x3x4x6_subscript0_share1       , x2x3x5x6_subscript0_share1       , x2x5x6x7_subscript0_share1       , x4x5x6x7_subscript0_share1       , x0x1x2x4_subscript0_share1       , x0x1x6x7_subscript0_share1       , x0x2x6x7_subscript0_share1       , x0x3x6x7_subscript0_share1       , x0x5x6x7_subscript0_share1       , x1x2x4x5_subscript0_share1       , x0x1x3x7_subscript0_share1       , x0x1x5x7_subscript0_share1       , x0x1x2x3x4_subscript0_share1     , x0x1x2x3x6_subscript0_share1     , x0x1x2x3x7_subscript0_share1     , x0x1x2x4x5_subscript0_share1     , x0x1x2x4x7_subscript0_share1     , x0x1x2x5x7_subscript0_share1     , x0x1x2x6x7_subscript0_share1     , x0x1x3x4x6_subscript0_share1     , x0x1x3x5x6_subscript0_share1     , x0x1x3x5x7_subscript0_share1     , x0x1x3x6x7_subscript0_share1     , x0x1x4x5x6_subscript0_share1     , x0x1x5x6x7_subscript0_share1     , x0x2x3x4x5_subscript0_share1     , x0x2x3x4x6_subscript0_share1     , x0x2x4x5x7_subscript0_share1     , x0x2x4x6x7_subscript0_share1     , x0x3x4x5x6_subscript0_share1     , x0x3x4x5x7_subscript0_share1     , x0x3x4x6x7_subscript0_share1     , x0x3x5x6x7_subscript0_share1     , x1x2x3x5x6_subscript0_share1     , x1x2x3x5x7_subscript0_share1     , x1x2x4x5x6_subscript0_share1     , x1x2x4x6x7_subscript0_share1     , x1x2x5x6x7_subscript0_share1     , x1x3x4x5x7_subscript0_share1     , x2x3x4x5x6_subscript0_share1     , x2x3x4x5x7_subscript0_share1     , x2x4x5x6x7_subscript0_share1     , x0x1x2x4x6_subscript0_share1     , x0x1x3x4x7_subscript0_share1     , x0x2x3x4x7_subscript0_share1     , x0x2x3x5x7_subscript0_share1     , x0x2x3x6x7_subscript0_share1     , x0x2x4x5x6_subscript0_share1     , x0x2x5x6x7_subscript0_share1     , x0x4x5x6x7_subscript0_share1     , x1x2x3x4x6_subscript0_share1     , x1x3x4x5x6_subscript0_share1     , x2x3x4x6x7_subscript0_share1     , x0x1x2x3x5_subscript0_share1     , x0x1x4x6x7_subscript0_share1     , x1x2x3x4x5_subscript0_share1     , x1x2x3x6x7_subscript0_share1     , x1x2x4x5x7_subscript0_share1     , x1x3x4x6x7_subscript0_share1     , x1x3x5x6x7_subscript0_share1     , x1x4x5x6x7_subscript0_share1     , x2x3x5x6x7_subscript0_share1     , x3x4x5x6x7_subscript0_share1     , x0x1x2x5x6_subscript0_share1     , x0x1x3x4x5_subscript0_share1     , x0x1x4x5x7_subscript0_share1     , x0x2x3x5x6_subscript0_share1     , x1x2x3x4x7_subscript0_share1     , x0x1x2x3x4x6_subscript0_share1   , x0x1x2x3x4x7_subscript0_share1   , x0x1x2x3x5x7_subscript0_share1   , x0x1x2x3x6x7_subscript0_share1   , x0x1x2x4x5x7_subscript0_share1   , x0x1x2x5x6x7_subscript0_share1   , x0x1x3x4x6x7_subscript0_share1   , x0x1x4x5x6x7_subscript0_share1   , x0x2x3x4x5x6_subscript0_share1   , x0x2x3x4x5x7_subscript0_share1   , x0x2x3x5x6x7_subscript0_share1   , x1x2x3x4x6x7_subscript0_share1   , x1x2x4x5x6x7_subscript0_share1   , x1x3x4x5x6x7_subscript0_share1   , x2x3x4x5x6x7_subscript0_share1   , x0x1x2x3x5x6_subscript0_share1   , x0x1x2x4x6x7_subscript0_share1   , x0x1x3x4x5x6_subscript0_share1   , x0x2x3x4x6x7_subscript0_share1   , x1x2x3x4x5x6_subscript0_share1   , x1x2x3x5x6x7_subscript0_share1   , x0x1x2x3x4x5_subscript0_share1   , x0x1x2x4x5x6_subscript0_share1   , x0x1x3x4x5x7_subscript0_share1   , x0x1x3x5x6x7_subscript0_share1   , x0x2x4x5x6x7_subscript0_share1   , x1x2x3x4x5x7_subscript0_share1   , x0x3x4x5x6x7_subscript0_share1   , x0x1x2x3x4x6x7_subscript0_share1 , x0x1x2x4x5x6x7_subscript0_share1 , x0x2x3x4x5x6x7_subscript0_share1 , x0x1x2x3x5x6x7_subscript0_share1 , x0x1x3x4x5x6x7_subscript0_share1 , x1x2x3x4x5x6x7_subscript0_share1 , x0x1x2x3x4x5x6_subscript0_share1 , x0x1x2x3x4x5x7_subscript0_share1
);

// Register stage

register_array_AES_oneshare first_cycle_share1_reg (
        clk,
        x0_subscript0_share1             , x1_subscript0_share1             , x2_subscript0_share1             , x3_subscript0_share1             , x4_subscript0_share1             , x5_subscript0_share1             , x6_subscript0_share1             , x7_subscript0_share1             , x0x1_subscript0_share1           , x0x4_subscript0_share1           , x0x5_subscript0_share1           , x0x6_subscript0_share1           , x1x2_subscript0_share1           , x1x3_subscript0_share1           , x1x4_subscript0_share1           , x1x6_subscript0_share1           , x2x3_subscript0_share1           , x2x4_subscript0_share1           , x2x6_subscript0_share1           , x2x7_subscript0_share1           , x4x6_subscript0_share1           , x5x6_subscript0_share1           , x5x7_subscript0_share1           , x6x7_subscript0_share1           , x0x2_subscript0_share1           , x0x3_subscript0_share1           , x0x7_subscript0_share1           , x1x7_subscript0_share1           , x3x7_subscript0_share1           , x4x5_subscript0_share1           , x3x4_subscript0_share1           , x4x7_subscript0_share1           , x3x6_subscript0_share1           , x1x5_subscript0_share1           , x2x5_subscript0_share1           , x3x5_subscript0_share1           , x0x1x4_subscript0_share1         , x0x1x6_subscript0_share1         , x0x1x7_subscript0_share1         , x0x2x4_subscript0_share1         , x0x2x5_subscript0_share1         , x0x2x6_subscript0_share1         , x0x2x7_subscript0_share1         , x0x3x4_subscript0_share1         , x0x3x5_subscript0_share1         , x0x3x6_subscript0_share1         , x0x4x6_subscript0_share1         , x0x4x7_subscript0_share1         , x1x2x3_subscript0_share1         , x1x2x4_subscript0_share1         , x1x2x6_subscript0_share1         , x1x3x4_subscript0_share1         , x1x3x7_subscript0_share1         , x1x4x6_subscript0_share1         , x1x5x6_subscript0_share1         , x2x3x5_subscript0_share1         , x2x3x7_subscript0_share1         , x2x4x7_subscript0_share1         , x2x5x6_subscript0_share1         , x2x5x7_subscript0_share1         , x2x6x7_subscript0_share1         , x3x4x7_subscript0_share1         , x3x5x7_subscript0_share1         , x3x6x7_subscript0_share1         , x4x5x6_subscript0_share1         , x5x6x7_subscript0_share1         , x0x1x3_subscript0_share1         , x0x2x3_subscript0_share1         , x0x4x5_subscript0_share1         , x0x5x7_subscript0_share1         , x0x6x7_subscript0_share1         , x1x3x5_subscript0_share1         , x1x3x6_subscript0_share1         , x1x4x7_subscript0_share1         , x2x3x4_subscript0_share1         , x2x3x6_subscript0_share1         , x3x4x6_subscript0_share1         , x3x5x6_subscript0_share1         , x0x1x5_subscript0_share1         , x0x3x7_subscript0_share1         , x1x2x5_subscript0_share1         , x1x2x7_subscript0_share1         , x1x4x5_subscript0_share1         , x1x5x7_subscript0_share1         , x2x4x5_subscript0_share1         , x3x4x5_subscript0_share1         , x4x6x7_subscript0_share1         , x1x6x7_subscript0_share1         , x4x5x7_subscript0_share1         , x0x1x2_subscript0_share1         , x0x5x6_subscript0_share1         , x2x4x6_subscript0_share1         , x0x1x2x3_subscript0_share1       , x0x1x2x5_subscript0_share1       , x0x1x2x6_subscript0_share1       , x0x1x2x7_subscript0_share1       , x0x1x4x5_subscript0_share1       , x0x1x4x7_subscript0_share1       , x0x2x3x5_subscript0_share1       , x0x2x3x7_subscript0_share1       , x0x2x4x5_subscript0_share1       , x0x2x4x7_subscript0_share1       , x0x2x5x6_subscript0_share1       , x0x2x5x7_subscript0_share1       , x0x3x4x6_subscript0_share1       , x0x3x5x6_subscript0_share1       , x0x4x5x6_subscript0_share1       , x0x4x5x7_subscript0_share1       , x0x4x6x7_subscript0_share1       , x1x2x3x5_subscript0_share1       , x1x2x3x6_subscript0_share1       , x1x2x3x7_subscript0_share1       , x1x2x4x6_subscript0_share1       , x1x2x4x7_subscript0_share1       , x1x2x6x7_subscript0_share1       , x1x3x4x6_subscript0_share1       , x1x3x6x7_subscript0_share1       , x1x4x5x6_subscript0_share1       , x1x4x5x7_subscript0_share1       , x1x5x6x7_subscript0_share1       , x2x3x5x7_subscript0_share1       , x2x3x6x7_subscript0_share1       , x2x4x5x6_subscript0_share1       , x2x4x5x7_subscript0_share1       , x3x5x6x7_subscript0_share1       , x0x1x3x4_subscript0_share1       , x0x1x3x6_subscript0_share1       , x0x1x5x6_subscript0_share1       , x0x2x3x6_subscript0_share1       , x0x3x4x5_subscript0_share1       , x1x2x5x6_subscript0_share1       , x1x2x5x7_subscript0_share1       , x1x3x4x5_subscript0_share1       , x1x3x4x7_subscript0_share1       , x1x3x5x6_subscript0_share1       , x1x3x5x7_subscript0_share1       , x1x4x6x7_subscript0_share1       , x2x3x4x5_subscript0_share1       , x2x3x4x7_subscript0_share1       , x2x4x6x7_subscript0_share1       , x3x4x5x6_subscript0_share1       , x3x4x5x7_subscript0_share1       , x3x4x6x7_subscript0_share1       , x0x1x3x5_subscript0_share1       , x0x1x4x6_subscript0_share1       , x0x2x3x4_subscript0_share1       , x0x2x4x6_subscript0_share1       , x0x3x4x7_subscript0_share1       , x0x3x5x7_subscript0_share1       , x1x2x3x4_subscript0_share1       , x2x3x4x6_subscript0_share1       , x2x3x5x6_subscript0_share1       , x2x5x6x7_subscript0_share1       , x4x5x6x7_subscript0_share1       , x0x1x2x4_subscript0_share1       , x0x1x6x7_subscript0_share1       , x0x2x6x7_subscript0_share1       , x0x3x6x7_subscript0_share1       , x0x5x6x7_subscript0_share1       , x1x2x4x5_subscript0_share1       , x0x1x3x7_subscript0_share1       , x0x1x5x7_subscript0_share1       , x0x1x2x3x4_subscript0_share1     , x0x1x2x3x6_subscript0_share1     , x0x1x2x3x7_subscript0_share1     , x0x1x2x4x5_subscript0_share1     , x0x1x2x4x7_subscript0_share1     , x0x1x2x5x7_subscript0_share1     , x0x1x2x6x7_subscript0_share1     , x0x1x3x4x6_subscript0_share1     , x0x1x3x5x6_subscript0_share1     , x0x1x3x5x7_subscript0_share1     , x0x1x3x6x7_subscript0_share1     , x0x1x4x5x6_subscript0_share1     , x0x1x5x6x7_subscript0_share1     , x0x2x3x4x5_subscript0_share1     , x0x2x3x4x6_subscript0_share1     , x0x2x4x5x7_subscript0_share1     , x0x2x4x6x7_subscript0_share1     , x0x3x4x5x6_subscript0_share1     , x0x3x4x5x7_subscript0_share1     , x0x3x4x6x7_subscript0_share1     , x0x3x5x6x7_subscript0_share1     , x1x2x3x5x6_subscript0_share1     , x1x2x3x5x7_subscript0_share1     , x1x2x4x5x6_subscript0_share1     , x1x2x4x6x7_subscript0_share1     , x1x2x5x6x7_subscript0_share1     , x1x3x4x5x7_subscript0_share1     , x2x3x4x5x6_subscript0_share1     , x2x3x4x5x7_subscript0_share1     , x2x4x5x6x7_subscript0_share1     , x0x1x2x4x6_subscript0_share1     , x0x1x3x4x7_subscript0_share1     , x0x2x3x4x7_subscript0_share1     , x0x2x3x5x7_subscript0_share1     , x0x2x3x6x7_subscript0_share1     , x0x2x4x5x6_subscript0_share1     , x0x2x5x6x7_subscript0_share1     , x0x4x5x6x7_subscript0_share1     , x1x2x3x4x6_subscript0_share1     , x1x3x4x5x6_subscript0_share1     , x2x3x4x6x7_subscript0_share1     , x0x1x2x3x5_subscript0_share1     , x0x1x4x6x7_subscript0_share1     , x1x2x3x4x5_subscript0_share1     , x1x2x3x6x7_subscript0_share1     , x1x2x4x5x7_subscript0_share1     , x1x3x4x6x7_subscript0_share1     , x1x3x5x6x7_subscript0_share1     , x1x4x5x6x7_subscript0_share1     , x2x3x5x6x7_subscript0_share1     , x3x4x5x6x7_subscript0_share1     , x0x1x2x5x6_subscript0_share1     , x0x1x3x4x5_subscript0_share1     , x0x1x4x5x7_subscript0_share1     , x0x2x3x5x6_subscript0_share1     , x1x2x3x4x7_subscript0_share1     , x0x1x2x3x4x6_subscript0_share1   , x0x1x2x3x4x7_subscript0_share1   , x0x1x2x3x5x7_subscript0_share1   , x0x1x2x3x6x7_subscript0_share1   , x0x1x2x4x5x7_subscript0_share1   , x0x1x2x5x6x7_subscript0_share1   , x0x1x3x4x6x7_subscript0_share1   , x0x1x4x5x6x7_subscript0_share1   , x0x2x3x4x5x6_subscript0_share1   , x0x2x3x4x5x7_subscript0_share1   , x0x2x3x5x6x7_subscript0_share1   , x1x2x3x4x6x7_subscript0_share1   , x1x2x4x5x6x7_subscript0_share1   , x1x3x4x5x6x7_subscript0_share1   , x2x3x4x5x6x7_subscript0_share1   , x0x1x2x3x5x6_subscript0_share1   , x0x1x2x4x6x7_subscript0_share1   , x0x1x3x4x5x6_subscript0_share1   , x0x2x3x4x6x7_subscript0_share1   , x1x2x3x4x5x6_subscript0_share1   , x1x2x3x5x6x7_subscript0_share1   , x0x1x2x3x4x5_subscript0_share1   , x0x1x2x4x5x6_subscript0_share1   , x0x1x3x4x5x7_subscript0_share1   , x0x1x3x5x6x7_subscript0_share1   , x0x2x4x5x6x7_subscript0_share1   , x1x2x3x4x5x7_subscript0_share1   , x0x3x4x5x6x7_subscript0_share1   , x0x1x2x3x4x6x7_subscript0_share1 , x0x1x2x4x5x6x7_subscript0_share1 , x0x2x3x4x5x6x7_subscript0_share1 , x0x1x2x3x5x6x7_subscript0_share1 , x0x1x3x4x5x6x7_subscript0_share1 , x1x2x3x4x5x6x7_subscript0_share1 , x0x1x2x3x4x5x6_subscript0_share1 , x0x1x2x3x4x5x7_subscript0_share1 ,
        x0_subscript0_share1_reg             , x1_subscript0_share1_reg             , x2_subscript0_share1_reg             , x3_subscript0_share1_reg             , x4_subscript0_share1_reg             , x5_subscript0_share1_reg             , x6_subscript0_share1_reg             , x7_subscript0_share1_reg             , x0x1_subscript0_share1_reg           , x0x4_subscript0_share1_reg           , x0x5_subscript0_share1_reg           , x0x6_subscript0_share1_reg           , x1x2_subscript0_share1_reg           , x1x3_subscript0_share1_reg           , x1x4_subscript0_share1_reg           , x1x6_subscript0_share1_reg           , x2x3_subscript0_share1_reg           , x2x4_subscript0_share1_reg           , x2x6_subscript0_share1_reg           , x2x7_subscript0_share1_reg           , x4x6_subscript0_share1_reg           , x5x6_subscript0_share1_reg           , x5x7_subscript0_share1_reg           , x6x7_subscript0_share1_reg           , x0x2_subscript0_share1_reg           , x0x3_subscript0_share1_reg           , x0x7_subscript0_share1_reg           , x1x7_subscript0_share1_reg           , x3x7_subscript0_share1_reg           , x4x5_subscript0_share1_reg           , x3x4_subscript0_share1_reg           , x4x7_subscript0_share1_reg           , x3x6_subscript0_share1_reg           , x1x5_subscript0_share1_reg           , x2x5_subscript0_share1_reg           , x3x5_subscript0_share1_reg           , x0x1x4_subscript0_share1_reg         , x0x1x6_subscript0_share1_reg         , x0x1x7_subscript0_share1_reg         , x0x2x4_subscript0_share1_reg         , x0x2x5_subscript0_share1_reg         , x0x2x6_subscript0_share1_reg         , x0x2x7_subscript0_share1_reg         , x0x3x4_subscript0_share1_reg         , x0x3x5_subscript0_share1_reg         , x0x3x6_subscript0_share1_reg         , x0x4x6_subscript0_share1_reg         , x0x4x7_subscript0_share1_reg         , x1x2x3_subscript0_share1_reg         , x1x2x4_subscript0_share1_reg         , x1x2x6_subscript0_share1_reg         , x1x3x4_subscript0_share1_reg         , x1x3x7_subscript0_share1_reg         , x1x4x6_subscript0_share1_reg         , x1x5x6_subscript0_share1_reg         , x2x3x5_subscript0_share1_reg         , x2x3x7_subscript0_share1_reg         , x2x4x7_subscript0_share1_reg         , x2x5x6_subscript0_share1_reg         , x2x5x7_subscript0_share1_reg         , x2x6x7_subscript0_share1_reg         , x3x4x7_subscript0_share1_reg         , x3x5x7_subscript0_share1_reg         , x3x6x7_subscript0_share1_reg         , x4x5x6_subscript0_share1_reg         , x5x6x7_subscript0_share1_reg         , x0x1x3_subscript0_share1_reg         , x0x2x3_subscript0_share1_reg         , x0x4x5_subscript0_share1_reg         , x0x5x7_subscript0_share1_reg         , x0x6x7_subscript0_share1_reg         , x1x3x5_subscript0_share1_reg         , x1x3x6_subscript0_share1_reg         , x1x4x7_subscript0_share1_reg         , x2x3x4_subscript0_share1_reg         , x2x3x6_subscript0_share1_reg         , x3x4x6_subscript0_share1_reg         , x3x5x6_subscript0_share1_reg         , x0x1x5_subscript0_share1_reg         , x0x3x7_subscript0_share1_reg         , x1x2x5_subscript0_share1_reg         , x1x2x7_subscript0_share1_reg         , x1x4x5_subscript0_share1_reg         , x1x5x7_subscript0_share1_reg         , x2x4x5_subscript0_share1_reg         , x3x4x5_subscript0_share1_reg         , x4x6x7_subscript0_share1_reg         , x1x6x7_subscript0_share1_reg         , x4x5x7_subscript0_share1_reg         , x0x1x2_subscript0_share1_reg         , x0x5x6_subscript0_share1_reg         , x2x4x6_subscript0_share1_reg         , x0x1x2x3_subscript0_share1_reg       , x0x1x2x5_subscript0_share1_reg       , x0x1x2x6_subscript0_share1_reg       , x0x1x2x7_subscript0_share1_reg       , x0x1x4x5_subscript0_share1_reg       , x0x1x4x7_subscript0_share1_reg       , x0x2x3x5_subscript0_share1_reg       , x0x2x3x7_subscript0_share1_reg       , x0x2x4x5_subscript0_share1_reg       , x0x2x4x7_subscript0_share1_reg       , x0x2x5x6_subscript0_share1_reg       , x0x2x5x7_subscript0_share1_reg       , x0x3x4x6_subscript0_share1_reg       , x0x3x5x6_subscript0_share1_reg       , x0x4x5x6_subscript0_share1_reg       , x0x4x5x7_subscript0_share1_reg       , x0x4x6x7_subscript0_share1_reg       , x1x2x3x5_subscript0_share1_reg       , x1x2x3x6_subscript0_share1_reg       , x1x2x3x7_subscript0_share1_reg       , x1x2x4x6_subscript0_share1_reg       , x1x2x4x7_subscript0_share1_reg       , x1x2x6x7_subscript0_share1_reg       , x1x3x4x6_subscript0_share1_reg       , x1x3x6x7_subscript0_share1_reg       , x1x4x5x6_subscript0_share1_reg       , x1x4x5x7_subscript0_share1_reg       , x1x5x6x7_subscript0_share1_reg       , x2x3x5x7_subscript0_share1_reg       , x2x3x6x7_subscript0_share1_reg       , x2x4x5x6_subscript0_share1_reg       , x2x4x5x7_subscript0_share1_reg       , x3x5x6x7_subscript0_share1_reg       , x0x1x3x4_subscript0_share1_reg       , x0x1x3x6_subscript0_share1_reg       , x0x1x5x6_subscript0_share1_reg       , x0x2x3x6_subscript0_share1_reg       , x0x3x4x5_subscript0_share1_reg       , x1x2x5x6_subscript0_share1_reg       , x1x2x5x7_subscript0_share1_reg       , x1x3x4x5_subscript0_share1_reg       , x1x3x4x7_subscript0_share1_reg       , x1x3x5x6_subscript0_share1_reg       , x1x3x5x7_subscript0_share1_reg       , x1x4x6x7_subscript0_share1_reg       , x2x3x4x5_subscript0_share1_reg       , x2x3x4x7_subscript0_share1_reg       , x2x4x6x7_subscript0_share1_reg       , x3x4x5x6_subscript0_share1_reg       , x3x4x5x7_subscript0_share1_reg       , x3x4x6x7_subscript0_share1_reg       , x0x1x3x5_subscript0_share1_reg       , x0x1x4x6_subscript0_share1_reg       , x0x2x3x4_subscript0_share1_reg       , x0x2x4x6_subscript0_share1_reg       , x0x3x4x7_subscript0_share1_reg       , x0x3x5x7_subscript0_share1_reg       , x1x2x3x4_subscript0_share1_reg       , x2x3x4x6_subscript0_share1_reg       , x2x3x5x6_subscript0_share1_reg       , x2x5x6x7_subscript0_share1_reg       , x4x5x6x7_subscript0_share1_reg       , x0x1x2x4_subscript0_share1_reg       , x0x1x6x7_subscript0_share1_reg       , x0x2x6x7_subscript0_share1_reg       , x0x3x6x7_subscript0_share1_reg       , x0x5x6x7_subscript0_share1_reg       , x1x2x4x5_subscript0_share1_reg       , x0x1x3x7_subscript0_share1_reg       , x0x1x5x7_subscript0_share1_reg       , x0x1x2x3x4_subscript0_share1_reg     , x0x1x2x3x6_subscript0_share1_reg     , x0x1x2x3x7_subscript0_share1_reg     , x0x1x2x4x5_subscript0_share1_reg     , x0x1x2x4x7_subscript0_share1_reg     , x0x1x2x5x7_subscript0_share1_reg     , x0x1x2x6x7_subscript0_share1_reg     , x0x1x3x4x6_subscript0_share1_reg     , x0x1x3x5x6_subscript0_share1_reg     , x0x1x3x5x7_subscript0_share1_reg     , x0x1x3x6x7_subscript0_share1_reg     , x0x1x4x5x6_subscript0_share1_reg     , x0x1x5x6x7_subscript0_share1_reg     , x0x2x3x4x5_subscript0_share1_reg     , x0x2x3x4x6_subscript0_share1_reg     , x0x2x4x5x7_subscript0_share1_reg     , x0x2x4x6x7_subscript0_share1_reg     , x0x3x4x5x6_subscript0_share1_reg     , x0x3x4x5x7_subscript0_share1_reg     , x0x3x4x6x7_subscript0_share1_reg     , x0x3x5x6x7_subscript0_share1_reg     , x1x2x3x5x6_subscript0_share1_reg     , x1x2x3x5x7_subscript0_share1_reg     , x1x2x4x5x6_subscript0_share1_reg     , x1x2x4x6x7_subscript0_share1_reg     , x1x2x5x6x7_subscript0_share1_reg     , x1x3x4x5x7_subscript0_share1_reg     , x2x3x4x5x6_subscript0_share1_reg     , x2x3x4x5x7_subscript0_share1_reg     , x2x4x5x6x7_subscript0_share1_reg     , x0x1x2x4x6_subscript0_share1_reg     , x0x1x3x4x7_subscript0_share1_reg     , x0x2x3x4x7_subscript0_share1_reg     , x0x2x3x5x7_subscript0_share1_reg     , x0x2x3x6x7_subscript0_share1_reg     , x0x2x4x5x6_subscript0_share1_reg     , x0x2x5x6x7_subscript0_share1_reg     , x0x4x5x6x7_subscript0_share1_reg     , x1x2x3x4x6_subscript0_share1_reg     , x1x3x4x5x6_subscript0_share1_reg     , x2x3x4x6x7_subscript0_share1_reg     , x0x1x2x3x5_subscript0_share1_reg     , x0x1x4x6x7_subscript0_share1_reg     , x1x2x3x4x5_subscript0_share1_reg     , x1x2x3x6x7_subscript0_share1_reg     , x1x2x4x5x7_subscript0_share1_reg     , x1x3x4x6x7_subscript0_share1_reg     , x1x3x5x6x7_subscript0_share1_reg     , x1x4x5x6x7_subscript0_share1_reg     , x2x3x5x6x7_subscript0_share1_reg     , x3x4x5x6x7_subscript0_share1_reg     , x0x1x2x5x6_subscript0_share1_reg     , x0x1x3x4x5_subscript0_share1_reg     , x0x1x4x5x7_subscript0_share1_reg     , x0x2x3x5x6_subscript0_share1_reg     , x1x2x3x4x7_subscript0_share1_reg     , x0x1x2x3x4x6_subscript0_share1_reg   , x0x1x2x3x4x7_subscript0_share1_reg   , x0x1x2x3x5x7_subscript0_share1_reg   , x0x1x2x3x6x7_subscript0_share1_reg   , x0x1x2x4x5x7_subscript0_share1_reg   , x0x1x2x5x6x7_subscript0_share1_reg   , x0x1x3x4x6x7_subscript0_share1_reg   , x0x1x4x5x6x7_subscript0_share1_reg   , x0x2x3x4x5x6_subscript0_share1_reg   , x0x2x3x4x5x7_subscript0_share1_reg   , x0x2x3x5x6x7_subscript0_share1_reg   , x1x2x3x4x6x7_subscript0_share1_reg   , x1x2x4x5x6x7_subscript0_share1_reg   , x1x3x4x5x6x7_subscript0_share1_reg   , x2x3x4x5x6x7_subscript0_share1_reg   , x0x1x2x3x5x6_subscript0_share1_reg   , x0x1x2x4x6x7_subscript0_share1_reg   , x0x1x3x4x5x6_subscript0_share1_reg   , x0x2x3x4x6x7_subscript0_share1_reg   , x1x2x3x4x5x6_subscript0_share1_reg   , x1x2x3x5x6x7_subscript0_share1_reg   , x0x1x2x3x4x5_subscript0_share1_reg   , x0x1x2x4x5x6_subscript0_share1_reg   , x0x1x3x4x5x7_subscript0_share1_reg   , x0x1x3x5x6x7_subscript0_share1_reg   , x0x2x4x5x6x7_subscript0_share1_reg   , x1x2x3x4x5x7_subscript0_share1_reg   , x0x3x4x5x6x7_subscript0_share1_reg   , x0x1x2x3x4x6x7_subscript0_share1_reg , x0x1x2x4x5x6x7_subscript0_share1_reg , x0x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x5x6x7_subscript0_share1_reg , x0x1x3x4x5x6x7_subscript0_share1_reg , x1x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x4x5x6_subscript0_share1_reg , x0x1x2x3x4x5x7_subscript0_share1_reg 
);
register_array_AES_oneshare first_cycle_share2_reg (
        clk,
        rand_first_cycle[1] ,rand_first_cycle[2] ,rand_first_cycle[3] ,rand_first_cycle[4] ,rand_first_cycle[5] ,rand_first_cycle[6] ,rand_first_cycle[7] ,rand_first_cycle[8] ,rand_first_cycle[9] ,rand_first_cycle[10] ,rand_first_cycle[11] ,rand_first_cycle[12] ,rand_first_cycle[13] ,rand_first_cycle[14] ,rand_first_cycle[15] ,rand_first_cycle[16] ,rand_first_cycle[17] ,rand_first_cycle[18] ,rand_first_cycle[19] ,rand_first_cycle[20] ,rand_first_cycle[21] ,rand_first_cycle[22] ,rand_first_cycle[23] ,rand_first_cycle[24] ,rand_first_cycle[25] ,rand_first_cycle[26] ,rand_first_cycle[27] ,rand_first_cycle[28] ,rand_first_cycle[29] ,rand_first_cycle[30] ,rand_first_cycle[31] ,rand_first_cycle[32] ,rand_first_cycle[33] ,rand_first_cycle[34] ,rand_first_cycle[35] ,rand_first_cycle[36] ,rand_first_cycle[37] ,rand_first_cycle[38] ,rand_first_cycle[39] ,rand_first_cycle[40] ,rand_first_cycle[41] ,rand_first_cycle[42] ,rand_first_cycle[43] ,rand_first_cycle[44] ,rand_first_cycle[45] ,rand_first_cycle[46] ,rand_first_cycle[47] ,rand_first_cycle[48] ,rand_first_cycle[49] ,rand_first_cycle[50] ,rand_first_cycle[51] ,rand_first_cycle[52] ,rand_first_cycle[53] ,rand_first_cycle[54] ,rand_first_cycle[55] ,rand_first_cycle[56] ,rand_first_cycle[57] ,rand_first_cycle[58] ,rand_first_cycle[59] ,rand_first_cycle[60] ,rand_first_cycle[61] ,rand_first_cycle[62] ,rand_first_cycle[63] ,rand_first_cycle[64] ,rand_first_cycle[65] ,rand_first_cycle[66] ,rand_first_cycle[67] ,rand_first_cycle[68] ,rand_first_cycle[69] ,rand_first_cycle[70] ,rand_first_cycle[71] ,rand_first_cycle[72] ,rand_first_cycle[73] ,rand_first_cycle[74] ,rand_first_cycle[75] ,rand_first_cycle[76] ,rand_first_cycle[77] ,rand_first_cycle[78] ,rand_first_cycle[79] ,rand_first_cycle[80] ,rand_first_cycle[81] ,rand_first_cycle[82] ,rand_first_cycle[83] ,rand_first_cycle[84] ,rand_first_cycle[85] ,rand_first_cycle[86] ,rand_first_cycle[87] ,rand_first_cycle[88] ,rand_first_cycle[89] ,rand_first_cycle[90] ,rand_first_cycle[91] ,rand_first_cycle[92] ,rand_first_cycle[93] ,rand_first_cycle[94] ,rand_first_cycle[95] ,rand_first_cycle[96] ,rand_first_cycle[97] ,rand_first_cycle[98] ,rand_first_cycle[99] ,rand_first_cycle[100] ,rand_first_cycle[101] ,rand_first_cycle[102] ,rand_first_cycle[103] ,rand_first_cycle[104] ,rand_first_cycle[105] ,rand_first_cycle[106] ,rand_first_cycle[107] ,rand_first_cycle[108] ,rand_first_cycle[109] ,rand_first_cycle[110] ,rand_first_cycle[111] ,rand_first_cycle[112] ,rand_first_cycle[113] ,rand_first_cycle[114] ,rand_first_cycle[115] ,rand_first_cycle[116] ,rand_first_cycle[117] ,rand_first_cycle[118] ,rand_first_cycle[119] ,rand_first_cycle[120] ,rand_first_cycle[121] ,rand_first_cycle[122] ,rand_first_cycle[123] ,rand_first_cycle[124] ,rand_first_cycle[125] ,rand_first_cycle[126] ,rand_first_cycle[127] ,rand_first_cycle[128] ,rand_first_cycle[129] ,rand_first_cycle[130] ,rand_first_cycle[131] ,rand_first_cycle[132] ,rand_first_cycle[133] ,rand_first_cycle[134] ,rand_first_cycle[135] ,rand_first_cycle[136] ,rand_first_cycle[137] ,rand_first_cycle[138] ,rand_first_cycle[139] ,rand_first_cycle[140] ,rand_first_cycle[141] ,rand_first_cycle[142] ,rand_first_cycle[143] ,rand_first_cycle[144] ,rand_first_cycle[145] ,rand_first_cycle[146] ,rand_first_cycle[147] ,rand_first_cycle[148] ,rand_first_cycle[149] ,rand_first_cycle[150] ,rand_first_cycle[151] ,rand_first_cycle[152] ,rand_first_cycle[153] ,rand_first_cycle[154] ,rand_first_cycle[155] ,rand_first_cycle[156] ,rand_first_cycle[157] ,rand_first_cycle[158] ,rand_first_cycle[159] ,rand_first_cycle[160] ,rand_first_cycle[161] ,rand_first_cycle[162] ,rand_first_cycle[163] ,rand_first_cycle[164] ,rand_first_cycle[165] ,rand_first_cycle[166] ,rand_first_cycle[167] ,rand_first_cycle[168] ,rand_first_cycle[169] ,rand_first_cycle[170] ,rand_first_cycle[171] ,rand_first_cycle[172] ,rand_first_cycle[173] ,rand_first_cycle[174] ,rand_first_cycle[175] ,rand_first_cycle[176] ,rand_first_cycle[177] ,rand_first_cycle[178] ,rand_first_cycle[179] ,rand_first_cycle[180] ,rand_first_cycle[181] ,rand_first_cycle[182] ,rand_first_cycle[183] ,rand_first_cycle[184] ,rand_first_cycle[185] ,rand_first_cycle[186] ,rand_first_cycle[187] ,rand_first_cycle[188] ,rand_first_cycle[189] ,rand_first_cycle[190] ,rand_first_cycle[191] ,rand_first_cycle[192] ,rand_first_cycle[193] ,rand_first_cycle[194] ,rand_first_cycle[195] ,rand_first_cycle[196] ,rand_first_cycle[197] ,rand_first_cycle[198] ,rand_first_cycle[199] ,rand_first_cycle[200] ,rand_first_cycle[201] ,rand_first_cycle[202] ,rand_first_cycle[203] ,rand_first_cycle[204] ,rand_first_cycle[205] ,rand_first_cycle[206] ,rand_first_cycle[207] ,rand_first_cycle[208] ,rand_first_cycle[209] ,rand_first_cycle[210] ,rand_first_cycle[211] ,rand_first_cycle[212] ,rand_first_cycle[213] ,rand_first_cycle[214] ,rand_first_cycle[215] ,rand_first_cycle[216] ,rand_first_cycle[217] ,rand_first_cycle[218] ,rand_first_cycle[219] ,rand_first_cycle[220] ,rand_first_cycle[221] ,rand_first_cycle[222] ,rand_first_cycle[223] ,rand_first_cycle[224] ,rand_first_cycle[225] ,rand_first_cycle[226] ,rand_first_cycle[227] ,rand_first_cycle[228] ,rand_first_cycle[229] ,rand_first_cycle[230] ,rand_first_cycle[231] ,rand_first_cycle[232] ,rand_first_cycle[233] ,rand_first_cycle[234] ,rand_first_cycle[235] ,rand_first_cycle[236] ,rand_first_cycle[237] ,rand_first_cycle[238] ,rand_first_cycle[239] ,rand_first_cycle[240] ,rand_first_cycle[241] ,rand_first_cycle[242] ,rand_first_cycle[243] ,rand_first_cycle[244] ,rand_first_cycle[245] ,rand_first_cycle[246] ,rand_first_cycle[247] ,rand_first_cycle[248] ,rand_first_cycle[249] ,rand_first_cycle[250] ,rand_first_cycle[251] ,rand_first_cycle[252] ,rand_first_cycle[253] ,rand_first_cycle[254] ,
        x0_subscript0_share2_reg             , x1_subscript0_share2_reg             , x2_subscript0_share2_reg             , x3_subscript0_share2_reg             , x4_subscript0_share2_reg             , x5_subscript0_share2_reg             , x6_subscript0_share2_reg             , x7_subscript0_share2_reg             , x0x1_subscript0_share2_reg           , x0x4_subscript0_share2_reg           , x0x5_subscript0_share2_reg           , x0x6_subscript0_share2_reg           , x1x2_subscript0_share2_reg           , x1x3_subscript0_share2_reg           , x1x4_subscript0_share2_reg           , x1x6_subscript0_share2_reg           , x2x3_subscript0_share2_reg           , x2x4_subscript0_share2_reg           , x2x6_subscript0_share2_reg           , x2x7_subscript0_share2_reg           , x4x6_subscript0_share2_reg           , x5x6_subscript0_share2_reg           , x5x7_subscript0_share2_reg           , x6x7_subscript0_share2_reg           , x0x2_subscript0_share2_reg           , x0x3_subscript0_share2_reg           , x0x7_subscript0_share2_reg           , x1x7_subscript0_share2_reg           , x3x7_subscript0_share2_reg           , x4x5_subscript0_share2_reg           , x3x4_subscript0_share2_reg           , x4x7_subscript0_share2_reg           , x3x6_subscript0_share2_reg           , x1x5_subscript0_share2_reg           , x2x5_subscript0_share2_reg           , x3x5_subscript0_share2_reg           , x0x1x4_subscript0_share2_reg         , x0x1x6_subscript0_share2_reg         , x0x1x7_subscript0_share2_reg         , x0x2x4_subscript0_share2_reg         , x0x2x5_subscript0_share2_reg         , x0x2x6_subscript0_share2_reg         , x0x2x7_subscript0_share2_reg         , x0x3x4_subscript0_share2_reg         , x0x3x5_subscript0_share2_reg         , x0x3x6_subscript0_share2_reg         , x0x4x6_subscript0_share2_reg         , x0x4x7_subscript0_share2_reg         , x1x2x3_subscript0_share2_reg         , x1x2x4_subscript0_share2_reg         , x1x2x6_subscript0_share2_reg         , x1x3x4_subscript0_share2_reg         , x1x3x7_subscript0_share2_reg         , x1x4x6_subscript0_share2_reg         , x1x5x6_subscript0_share2_reg         , x2x3x5_subscript0_share2_reg         , x2x3x7_subscript0_share2_reg         , x2x4x7_subscript0_share2_reg         , x2x5x6_subscript0_share2_reg         , x2x5x7_subscript0_share2_reg         , x2x6x7_subscript0_share2_reg         , x3x4x7_subscript0_share2_reg         , x3x5x7_subscript0_share2_reg         , x3x6x7_subscript0_share2_reg         , x4x5x6_subscript0_share2_reg         , x5x6x7_subscript0_share2_reg         , x0x1x3_subscript0_share2_reg         , x0x2x3_subscript0_share2_reg         , x0x4x5_subscript0_share2_reg         , x0x5x7_subscript0_share2_reg         , x0x6x7_subscript0_share2_reg         , x1x3x5_subscript0_share2_reg         , x1x3x6_subscript0_share2_reg         , x1x4x7_subscript0_share2_reg         , x2x3x4_subscript0_share2_reg         , x2x3x6_subscript0_share2_reg         , x3x4x6_subscript0_share2_reg         , x3x5x6_subscript0_share2_reg         , x0x1x5_subscript0_share2_reg         , x0x3x7_subscript0_share2_reg         , x1x2x5_subscript0_share2_reg         , x1x2x7_subscript0_share2_reg         , x1x4x5_subscript0_share2_reg         , x1x5x7_subscript0_share2_reg         , x2x4x5_subscript0_share2_reg         , x3x4x5_subscript0_share2_reg         , x4x6x7_subscript0_share2_reg         , x1x6x7_subscript0_share2_reg         , x4x5x7_subscript0_share2_reg         , x0x1x2_subscript0_share2_reg         , x0x5x6_subscript0_share2_reg         , x2x4x6_subscript0_share2_reg         , x0x1x2x3_subscript0_share2_reg       , x0x1x2x5_subscript0_share2_reg       , x0x1x2x6_subscript0_share2_reg       , x0x1x2x7_subscript0_share2_reg       , x0x1x4x5_subscript0_share2_reg       , x0x1x4x7_subscript0_share2_reg       , x0x2x3x5_subscript0_share2_reg       , x0x2x3x7_subscript0_share2_reg       , x0x2x4x5_subscript0_share2_reg       , x0x2x4x7_subscript0_share2_reg       , x0x2x5x6_subscript0_share2_reg       , x0x2x5x7_subscript0_share2_reg       , x0x3x4x6_subscript0_share2_reg       , x0x3x5x6_subscript0_share2_reg       , x0x4x5x6_subscript0_share2_reg       , x0x4x5x7_subscript0_share2_reg       , x0x4x6x7_subscript0_share2_reg       , x1x2x3x5_subscript0_share2_reg       , x1x2x3x6_subscript0_share2_reg       , x1x2x3x7_subscript0_share2_reg       , x1x2x4x6_subscript0_share2_reg       , x1x2x4x7_subscript0_share2_reg       , x1x2x6x7_subscript0_share2_reg       , x1x3x4x6_subscript0_share2_reg       , x1x3x6x7_subscript0_share2_reg       , x1x4x5x6_subscript0_share2_reg       , x1x4x5x7_subscript0_share2_reg       , x1x5x6x7_subscript0_share2_reg       , x2x3x5x7_subscript0_share2_reg       , x2x3x6x7_subscript0_share2_reg       , x2x4x5x6_subscript0_share2_reg       , x2x4x5x7_subscript0_share2_reg       , x3x5x6x7_subscript0_share2_reg       , x0x1x3x4_subscript0_share2_reg       , x0x1x3x6_subscript0_share2_reg       , x0x1x5x6_subscript0_share2_reg       , x0x2x3x6_subscript0_share2_reg       , x0x3x4x5_subscript0_share2_reg       , x1x2x5x6_subscript0_share2_reg       , x1x2x5x7_subscript0_share2_reg       , x1x3x4x5_subscript0_share2_reg       , x1x3x4x7_subscript0_share2_reg       , x1x3x5x6_subscript0_share2_reg       , x1x3x5x7_subscript0_share2_reg       , x1x4x6x7_subscript0_share2_reg       , x2x3x4x5_subscript0_share2_reg       , x2x3x4x7_subscript0_share2_reg       , x2x4x6x7_subscript0_share2_reg       , x3x4x5x6_subscript0_share2_reg       , x3x4x5x7_subscript0_share2_reg       , x3x4x6x7_subscript0_share2_reg       , x0x1x3x5_subscript0_share2_reg       , x0x1x4x6_subscript0_share2_reg       , x0x2x3x4_subscript0_share2_reg       , x0x2x4x6_subscript0_share2_reg       , x0x3x4x7_subscript0_share2_reg       , x0x3x5x7_subscript0_share2_reg       , x1x2x3x4_subscript0_share2_reg       , x2x3x4x6_subscript0_share2_reg       , x2x3x5x6_subscript0_share2_reg       , x2x5x6x7_subscript0_share2_reg       , x4x5x6x7_subscript0_share2_reg       , x0x1x2x4_subscript0_share2_reg       , x0x1x6x7_subscript0_share2_reg       , x0x2x6x7_subscript0_share2_reg       , x0x3x6x7_subscript0_share2_reg       , x0x5x6x7_subscript0_share2_reg       , x1x2x4x5_subscript0_share2_reg       , x0x1x3x7_subscript0_share2_reg       , x0x1x5x7_subscript0_share2_reg       , x0x1x2x3x4_subscript0_share2_reg     , x0x1x2x3x6_subscript0_share2_reg     , x0x1x2x3x7_subscript0_share2_reg     , x0x1x2x4x5_subscript0_share2_reg     , x0x1x2x4x7_subscript0_share2_reg     , x0x1x2x5x7_subscript0_share2_reg     , x0x1x2x6x7_subscript0_share2_reg     , x0x1x3x4x6_subscript0_share2_reg     , x0x1x3x5x6_subscript0_share2_reg     , x0x1x3x5x7_subscript0_share2_reg     , x0x1x3x6x7_subscript0_share2_reg     , x0x1x4x5x6_subscript0_share2_reg     , x0x1x5x6x7_subscript0_share2_reg     , x0x2x3x4x5_subscript0_share2_reg     , x0x2x3x4x6_subscript0_share2_reg     , x0x2x4x5x7_subscript0_share2_reg     , x0x2x4x6x7_subscript0_share2_reg     , x0x3x4x5x6_subscript0_share2_reg     , x0x3x4x5x7_subscript0_share2_reg     , x0x3x4x6x7_subscript0_share2_reg     , x0x3x5x6x7_subscript0_share2_reg     , x1x2x3x5x6_subscript0_share2_reg     , x1x2x3x5x7_subscript0_share2_reg     , x1x2x4x5x6_subscript0_share2_reg     , x1x2x4x6x7_subscript0_share2_reg     , x1x2x5x6x7_subscript0_share2_reg     , x1x3x4x5x7_subscript0_share2_reg     , x2x3x4x5x6_subscript0_share2_reg     , x2x3x4x5x7_subscript0_share2_reg     , x2x4x5x6x7_subscript0_share2_reg     , x0x1x2x4x6_subscript0_share2_reg     , x0x1x3x4x7_subscript0_share2_reg     , x0x2x3x4x7_subscript0_share2_reg     , x0x2x3x5x7_subscript0_share2_reg     , x0x2x3x6x7_subscript0_share2_reg     , x0x2x4x5x6_subscript0_share2_reg     , x0x2x5x6x7_subscript0_share2_reg     , x0x4x5x6x7_subscript0_share2_reg     , x1x2x3x4x6_subscript0_share2_reg     , x1x3x4x5x6_subscript0_share2_reg     , x2x3x4x6x7_subscript0_share2_reg     , x0x1x2x3x5_subscript0_share2_reg     , x0x1x4x6x7_subscript0_share2_reg     , x1x2x3x4x5_subscript0_share2_reg     , x1x2x3x6x7_subscript0_share2_reg     , x1x2x4x5x7_subscript0_share2_reg     , x1x3x4x6x7_subscript0_share2_reg     , x1x3x5x6x7_subscript0_share2_reg     , x1x4x5x6x7_subscript0_share2_reg     , x2x3x5x6x7_subscript0_share2_reg     , x3x4x5x6x7_subscript0_share2_reg     , x0x1x2x5x6_subscript0_share2_reg     , x0x1x3x4x5_subscript0_share2_reg     , x0x1x4x5x7_subscript0_share2_reg     , x0x2x3x5x6_subscript0_share2_reg     , x1x2x3x4x7_subscript0_share2_reg     , x0x1x2x3x4x6_subscript0_share2_reg   , x0x1x2x3x4x7_subscript0_share2_reg   , x0x1x2x3x5x7_subscript0_share2_reg   , x0x1x2x3x6x7_subscript0_share2_reg   , x0x1x2x4x5x7_subscript0_share2_reg   , x0x1x2x5x6x7_subscript0_share2_reg   , x0x1x3x4x6x7_subscript0_share2_reg   , x0x1x4x5x6x7_subscript0_share2_reg   , x0x2x3x4x5x6_subscript0_share2_reg   , x0x2x3x4x5x7_subscript0_share2_reg   , x0x2x3x5x6x7_subscript0_share2_reg   , x1x2x3x4x6x7_subscript0_share2_reg   , x1x2x4x5x6x7_subscript0_share2_reg   , x1x3x4x5x6x7_subscript0_share2_reg   , x2x3x4x5x6x7_subscript0_share2_reg   , x0x1x2x3x5x6_subscript0_share2_reg   , x0x1x2x4x6x7_subscript0_share2_reg   , x0x1x3x4x5x6_subscript0_share2_reg   , x0x2x3x4x6x7_subscript0_share2_reg   , x1x2x3x4x5x6_subscript0_share2_reg   , x1x2x3x5x6x7_subscript0_share2_reg   , x0x1x2x3x4x5_subscript0_share2_reg   , x0x1x2x4x5x6_subscript0_share2_reg   , x0x1x3x4x5x7_subscript0_share2_reg   , x0x1x3x5x6x7_subscript0_share2_reg   , x0x2x4x5x6x7_subscript0_share2_reg   , x1x2x3x4x5x7_subscript0_share2_reg   , x0x3x4x5x6x7_subscript0_share2_reg   , x0x1x2x3x4x6x7_subscript0_share2_reg , x0x1x2x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6x7_subscript0_share2_reg , x0x1x3x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5x6_subscript0_share2_reg , x0x1x2x3x4x5x7_subscript0_share2_reg 
);
register_array_8bit_AES  reg_first_cycle_pipeline_share2 (clk , x0_input_share2, x1_input_share2, x2_input_share2, x3_input_share2, x4_input_share2, x5_input_share2, x6_input_share2, x7_input_share2, x0_pipelined_share2_reg, x1_pipelined_share2_reg, x2_pipelined_share2_reg, x3_pipelined_share2_reg, x4_pipelined_share2_reg, x5_pipelined_share2_reg, x6_pipelined_share2_reg, x7_pipelined_share2_reg );
register_array_8bit_AES  reg_first_cycle_pipeline_share3 (clk , x0_input_share3, x1_input_share3, x2_input_share3, x3_input_share3, x4_input_share3, x5_input_share3, x6_input_share3, x7_input_share3, x0_pipelined_share3_reg, x1_pipelined_share3_reg, x2_pipelined_share3_reg, x3_pipelined_share3_reg, x4_pipelined_share3_reg, x5_pipelined_share3_reg, x6_pipelined_share3_reg, x7_pipelined_share3_reg );

// Second Cycle Logic 

combi_logic_cycle2_output_share1 inst_second_cycle_share1(
    x0_subscript0_share1_reg , x2_subscript0_share1_reg , x3_subscript0_share1_reg , x4_subscript0_share1_reg , x6_subscript0_share1_reg , x7_subscript0_share1_reg , x1_subscript0_share1_reg , x5_subscript0_share1_reg , x0x1_subscript0_share1_reg , x0x4_subscript0_share1_reg , x0x5_subscript0_share1_reg , x0x6_subscript0_share1_reg , x1x2_subscript0_share1_reg , x1x3_subscript0_share1_reg , x1x4_subscript0_share1_reg , x1x6_subscript0_share1_reg , x2x3_subscript0_share1_reg , x2x4_subscript0_share1_reg , x2x6_subscript0_share1_reg , x2x7_subscript0_share1_reg , x4x6_subscript0_share1_reg , x5x6_subscript0_share1_reg , x5x7_subscript0_share1_reg , x6x7_subscript0_share1_reg , x0x2_subscript0_share1_reg , x0x3_subscript0_share1_reg , x0x7_subscript0_share1_reg , x1x7_subscript0_share1_reg , x3x7_subscript0_share1_reg , x4x5_subscript0_share1_reg , x3x4_subscript0_share1_reg , x4x7_subscript0_share1_reg , x3x6_subscript0_share1_reg , x1x5_subscript0_share1_reg , x2x5_subscript0_share1_reg , x3x5_subscript0_share1_reg , x0x1x4_subscript0_share1_reg , x0x1x6_subscript0_share1_reg , x0x1x7_subscript0_share1_reg , x0x2x4_subscript0_share1_reg , x0x2x5_subscript0_share1_reg , x0x2x6_subscript0_share1_reg , x0x2x7_subscript0_share1_reg , x0x3x4_subscript0_share1_reg , x0x3x5_subscript0_share1_reg , x0x3x6_subscript0_share1_reg , x0x4x6_subscript0_share1_reg , x0x4x7_subscript0_share1_reg , x1x2x3_subscript0_share1_reg , x1x2x4_subscript0_share1_reg , x1x2x6_subscript0_share1_reg , x1x3x4_subscript0_share1_reg , x1x3x7_subscript0_share1_reg , x1x4x6_subscript0_share1_reg , x1x5x6_subscript0_share1_reg , x2x3x5_subscript0_share1_reg , x2x3x7_subscript0_share1_reg , x2x4x7_subscript0_share1_reg , x2x5x6_subscript0_share1_reg , x2x5x7_subscript0_share1_reg , x2x6x7_subscript0_share1_reg , x3x4x7_subscript0_share1_reg , x3x5x7_subscript0_share1_reg , x3x6x7_subscript0_share1_reg , x4x5x6_subscript0_share1_reg , x5x6x7_subscript0_share1_reg , x0x1x3_subscript0_share1_reg , x0x2x3_subscript0_share1_reg , x0x4x5_subscript0_share1_reg , x0x5x7_subscript0_share1_reg , x0x6x7_subscript0_share1_reg , x1x3x5_subscript0_share1_reg , x1x3x6_subscript0_share1_reg , x1x4x7_subscript0_share1_reg , x2x3x4_subscript0_share1_reg , x2x3x6_subscript0_share1_reg , x3x4x6_subscript0_share1_reg , x3x5x6_subscript0_share1_reg , x0x1x5_subscript0_share1_reg , x0x3x7_subscript0_share1_reg , x1x2x5_subscript0_share1_reg , x1x2x7_subscript0_share1_reg , x1x4x5_subscript0_share1_reg , x1x5x7_subscript0_share1_reg , x2x4x5_subscript0_share1_reg , x3x4x5_subscript0_share1_reg , x4x6x7_subscript0_share1_reg , x1x6x7_subscript0_share1_reg , x4x5x7_subscript0_share1_reg , x0x1x2_subscript0_share1_reg , x0x5x6_subscript0_share1_reg , x2x4x6_subscript0_share1_reg , x0x1x2x3_subscript0_share1_reg , x0x1x2x5_subscript0_share1_reg , x0x1x2x6_subscript0_share1_reg , x0x1x2x7_subscript0_share1_reg , x0x1x4x5_subscript0_share1_reg , x0x1x4x7_subscript0_share1_reg , x0x2x3x5_subscript0_share1_reg , x0x2x3x7_subscript0_share1_reg , x0x2x4x5_subscript0_share1_reg , x0x2x4x7_subscript0_share1_reg , x0x2x5x6_subscript0_share1_reg , x0x2x5x7_subscript0_share1_reg , x0x3x4x6_subscript0_share1_reg , x0x3x5x6_subscript0_share1_reg , x0x4x5x6_subscript0_share1_reg , x0x4x5x7_subscript0_share1_reg , x0x4x6x7_subscript0_share1_reg , x1x2x3x5_subscript0_share1_reg , x1x2x3x6_subscript0_share1_reg , x1x2x3x7_subscript0_share1_reg , x1x2x4x6_subscript0_share1_reg , x1x2x4x7_subscript0_share1_reg , x1x2x6x7_subscript0_share1_reg , x1x3x4x6_subscript0_share1_reg , x1x3x6x7_subscript0_share1_reg , x1x4x5x6_subscript0_share1_reg , x1x4x5x7_subscript0_share1_reg , x1x5x6x7_subscript0_share1_reg , x2x3x5x7_subscript0_share1_reg , x2x3x6x7_subscript0_share1_reg , x2x4x5x6_subscript0_share1_reg , x2x4x5x7_subscript0_share1_reg , x3x5x6x7_subscript0_share1_reg , x0x1x3x4_subscript0_share1_reg , x0x1x3x6_subscript0_share1_reg , x0x1x5x6_subscript0_share1_reg , x0x2x3x6_subscript0_share1_reg , x0x3x4x5_subscript0_share1_reg , x1x2x5x6_subscript0_share1_reg , x1x2x5x7_subscript0_share1_reg , x1x3x4x5_subscript0_share1_reg , x1x3x4x7_subscript0_share1_reg , x1x3x5x6_subscript0_share1_reg , x1x3x5x7_subscript0_share1_reg , x1x4x6x7_subscript0_share1_reg , x2x3x4x5_subscript0_share1_reg , x2x3x4x7_subscript0_share1_reg , x2x4x6x7_subscript0_share1_reg , x3x4x5x6_subscript0_share1_reg , x3x4x5x7_subscript0_share1_reg , x3x4x6x7_subscript0_share1_reg , x0x1x3x5_subscript0_share1_reg , x0x1x4x6_subscript0_share1_reg , x0x2x3x4_subscript0_share1_reg , x0x2x4x6_subscript0_share1_reg , x0x3x4x7_subscript0_share1_reg , x0x3x5x7_subscript0_share1_reg , x1x2x3x4_subscript0_share1_reg , x2x3x4x6_subscript0_share1_reg , x2x3x5x6_subscript0_share1_reg , x2x5x6x7_subscript0_share1_reg , x4x5x6x7_subscript0_share1_reg , x0x1x2x4_subscript0_share1_reg , x0x1x6x7_subscript0_share1_reg , x0x2x6x7_subscript0_share1_reg , x0x3x6x7_subscript0_share1_reg , x0x5x6x7_subscript0_share1_reg , x1x2x4x5_subscript0_share1_reg , x0x1x3x7_subscript0_share1_reg , x0x1x5x7_subscript0_share1_reg , x0x1x2x3x4_subscript0_share1_reg , x0x1x2x3x6_subscript0_share1_reg , x0x1x2x3x7_subscript0_share1_reg , x0x1x2x4x5_subscript0_share1_reg , x0x1x2x4x7_subscript0_share1_reg , x0x1x2x5x7_subscript0_share1_reg , x0x1x2x6x7_subscript0_share1_reg , x0x1x3x4x6_subscript0_share1_reg , x0x1x3x5x6_subscript0_share1_reg , x0x1x3x5x7_subscript0_share1_reg , x0x1x3x6x7_subscript0_share1_reg , x0x1x4x5x6_subscript0_share1_reg , x0x1x5x6x7_subscript0_share1_reg , x0x2x3x4x5_subscript0_share1_reg , x0x2x3x4x6_subscript0_share1_reg , x0x2x4x5x7_subscript0_share1_reg , x0x2x4x6x7_subscript0_share1_reg , x0x3x4x5x6_subscript0_share1_reg , x0x3x4x5x7_subscript0_share1_reg , x0x3x4x6x7_subscript0_share1_reg , x0x3x5x6x7_subscript0_share1_reg , x1x2x3x5x6_subscript0_share1_reg , x1x2x3x5x7_subscript0_share1_reg , x1x2x4x5x6_subscript0_share1_reg , x1x2x4x6x7_subscript0_share1_reg , x1x2x5x6x7_subscript0_share1_reg , x1x3x4x5x7_subscript0_share1_reg , x2x3x4x5x6_subscript0_share1_reg , x2x3x4x5x7_subscript0_share1_reg , x2x4x5x6x7_subscript0_share1_reg , x0x1x2x4x6_subscript0_share1_reg , x0x1x3x4x7_subscript0_share1_reg , x0x2x3x4x7_subscript0_share1_reg , x0x2x3x5x7_subscript0_share1_reg , x0x2x3x6x7_subscript0_share1_reg , x0x2x4x5x6_subscript0_share1_reg , x0x2x5x6x7_subscript0_share1_reg , x0x4x5x6x7_subscript0_share1_reg , x1x2x3x4x6_subscript0_share1_reg , x1x3x4x5x6_subscript0_share1_reg , x2x3x4x6x7_subscript0_share1_reg , x0x1x2x3x5_subscript0_share1_reg , x0x1x4x6x7_subscript0_share1_reg , x1x2x3x4x5_subscript0_share1_reg , x1x2x3x6x7_subscript0_share1_reg , x1x2x4x5x7_subscript0_share1_reg , x1x3x4x6x7_subscript0_share1_reg , x1x3x5x6x7_subscript0_share1_reg , x1x4x5x6x7_subscript0_share1_reg , x2x3x5x6x7_subscript0_share1_reg , x3x4x5x6x7_subscript0_share1_reg , x0x1x2x5x6_subscript0_share1_reg , x0x1x3x4x5_subscript0_share1_reg , x0x1x4x5x7_subscript0_share1_reg , x0x2x3x5x6_subscript0_share1_reg , x1x2x3x4x7_subscript0_share1_reg , x0x1x2x3x4x6_subscript0_share1_reg , x0x1x2x3x4x7_subscript0_share1_reg , x0x1x2x3x5x7_subscript0_share1_reg , x0x1x2x3x6x7_subscript0_share1_reg , x0x1x2x4x5x7_subscript0_share1_reg , x0x1x2x5x6x7_subscript0_share1_reg , x0x1x3x4x6x7_subscript0_share1_reg , x0x1x4x5x6x7_subscript0_share1_reg , x0x2x3x4x5x6_subscript0_share1_reg , x0x2x3x4x5x7_subscript0_share1_reg , x0x2x3x5x6x7_subscript0_share1_reg , x1x2x3x4x6x7_subscript0_share1_reg , x1x2x4x5x6x7_subscript0_share1_reg , x1x3x4x5x6x7_subscript0_share1_reg , x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x5x6_subscript0_share1_reg , x0x1x2x4x6x7_subscript0_share1_reg , x0x1x3x4x5x6_subscript0_share1_reg , x0x2x3x4x6x7_subscript0_share1_reg , x1x2x3x4x5x6_subscript0_share1_reg , x1x2x3x5x6x7_subscript0_share1_reg , x0x1x2x3x4x5_subscript0_share1_reg , x0x1x2x4x5x6_subscript0_share1_reg , x0x1x3x4x5x7_subscript0_share1_reg , x0x1x3x5x6x7_subscript0_share1_reg , x0x2x4x5x6x7_subscript0_share1_reg , x1x2x3x4x5x7_subscript0_share1_reg , x0x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x4x6x7_subscript0_share1_reg , x0x1x2x4x5x6x7_subscript0_share1_reg , x0x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x5x6x7_subscript0_share1_reg , x0x1x3x4x5x6x7_subscript0_share1_reg , x1x2x3x4x5x6x7_subscript0_share1_reg , x0x1x2x3x4x5x6_subscript0_share1_reg , x0x1x2x3x4x5x7_subscript0_share1_reg , 
    x0_pipelined_share2_reg ,x1_pipelined_share2_reg ,x2_pipelined_share2_reg ,x3_pipelined_share2_reg ,x4_pipelined_share2_reg ,x5_pipelined_share2_reg ,x6_pipelined_share2_reg ,x7_pipelined_share2_reg ,
    x0_subscript1_share1, x1_subscript1_share1, x2_subscript1_share1, x3_subscript1_share1, x4_subscript1_share1, x5_subscript1_share1, x6_subscript1_share1, x7_subscript1_share1 , x0x1_subscript1_share1 , x0x2_subscript1_share1 , x0x3_subscript1_share1 , x0x4_subscript1_share1 , x0x5_subscript1_share1 , x0x6_subscript1_share1 , x0x7_subscript1_share1 , x1x2_subscript1_share1 , x1x3_subscript1_share1 , x1x4_subscript1_share1 , x1x5_subscript1_share1 , x1x6_subscript1_share1 , x1x7_subscript1_share1 , x2x3_subscript1_share1 , x2x4_subscript1_share1 , x2x5_subscript1_share1 , x2x6_subscript1_share1 , x2x7_subscript1_share1 , x3x4_subscript1_share1 , x3x5_subscript1_share1 , x3x6_subscript1_share1 , x3x7_subscript1_share1 , x4x5_subscript1_share1 , x4x6_subscript1_share1 , x4x7_subscript1_share1 , x5x6_subscript1_share1 , x5x7_subscript1_share1 , x6x7_subscript1_share1 , x0x1x2_subscript1_share1 , x0x1x3_subscript1_share1 , x0x1x4_subscript1_share1 , x0x1x5_subscript1_share1 , x0x1x6_subscript1_share1 , x0x1x7_subscript1_share1 , x0x2x3_subscript1_share1 , x0x2x4_subscript1_share1 , x0x2x5_subscript1_share1 , x0x2x6_subscript1_share1 , x0x2x7_subscript1_share1 , x0x3x4_subscript1_share1 , x0x3x5_subscript1_share1 , x0x3x6_subscript1_share1 , x0x3x7_subscript1_share1 , x0x4x5_subscript1_share1 , x0x4x6_subscript1_share1 , x0x4x7_subscript1_share1 , x0x5x6_subscript1_share1 , x0x5x7_subscript1_share1 , x0x6x7_subscript1_share1 , x1x2x3_subscript1_share1 , x1x2x4_subscript1_share1 , x1x2x5_subscript1_share1 , x1x2x6_subscript1_share1 , x1x2x7_subscript1_share1 , x1x3x4_subscript1_share1 , x1x3x5_subscript1_share1 , x1x3x6_subscript1_share1 , x1x3x7_subscript1_share1 , x1x4x5_subscript1_share1 , x1x4x6_subscript1_share1 , x1x4x7_subscript1_share1 , x1x5x6_subscript1_share1 , x1x5x7_subscript1_share1 , x1x6x7_subscript1_share1 , x2x3x4_subscript1_share1 , x2x3x5_subscript1_share1 , x2x3x6_subscript1_share1 , x2x3x7_subscript1_share1 , x2x4x5_subscript1_share1 , x2x4x6_subscript1_share1 , x2x4x7_subscript1_share1 , x2x5x6_subscript1_share1 , x2x5x7_subscript1_share1 , x2x6x7_subscript1_share1 , x3x4x5_subscript1_share1 , x3x4x6_subscript1_share1 , x3x4x7_subscript1_share1 , x3x5x6_subscript1_share1 , x3x5x7_subscript1_share1 , x3x6x7_subscript1_share1 , x4x5x6_subscript1_share1 , x4x5x7_subscript1_share1 , x4x6x7_subscript1_share1 , x5x6x7_subscript1_share1 , x0x1x2x3_subscript1_share1 , x0x1x2x4_subscript1_share1 , x0x1x2x5_subscript1_share1 , x0x1x2x6_subscript1_share1 , x0x1x2x7_subscript1_share1 , x0x1x3x4_subscript1_share1 , x0x1x3x5_subscript1_share1 , x0x1x3x6_subscript1_share1 , x0x1x3x7_subscript1_share1 , x0x1x4x5_subscript1_share1 , x0x1x4x6_subscript1_share1 , x0x1x4x7_subscript1_share1 , x0x1x5x6_subscript1_share1 , x0x1x5x7_subscript1_share1 , x0x1x6x7_subscript1_share1 , x0x2x3x4_subscript1_share1 , x0x2x3x5_subscript1_share1 , x0x2x3x6_subscript1_share1 , x0x2x3x7_subscript1_share1 , x0x2x4x5_subscript1_share1 , x0x2x4x6_subscript1_share1 , x0x2x4x7_subscript1_share1 , x0x2x5x6_subscript1_share1 , x0x2x5x7_subscript1_share1 , x0x2x6x7_subscript1_share1 , x0x3x4x5_subscript1_share1 , x0x3x4x6_subscript1_share1 , x0x3x4x7_subscript1_share1 , x0x3x5x6_subscript1_share1 , x0x3x5x7_subscript1_share1 , x0x3x6x7_subscript1_share1 , x0x4x5x6_subscript1_share1 , x0x4x5x7_subscript1_share1 , x0x4x6x7_subscript1_share1 , x0x5x6x7_subscript1_share1 , x1x2x3x4_subscript1_share1 , x1x2x3x5_subscript1_share1 , x1x2x3x6_subscript1_share1 , x1x2x3x7_subscript1_share1 , x1x2x4x5_subscript1_share1 , x1x2x4x6_subscript1_share1 , x1x2x4x7_subscript1_share1 , x1x2x5x6_subscript1_share1 , x1x2x5x7_subscript1_share1 , x1x2x6x7_subscript1_share1 , x1x3x4x5_subscript1_share1 , x1x3x4x6_subscript1_share1 , x1x3x4x7_subscript1_share1 , x1x3x5x6_subscript1_share1 , x1x3x5x7_subscript1_share1 , x1x3x6x7_subscript1_share1 , x1x4x5x6_subscript1_share1 , x1x4x5x7_subscript1_share1 , x1x4x6x7_subscript1_share1 , x1x5x6x7_subscript1_share1 , x2x3x4x5_subscript1_share1 , x2x3x4x6_subscript1_share1 , x2x3x4x7_subscript1_share1 , x2x3x5x6_subscript1_share1 , x2x3x5x7_subscript1_share1 , x2x3x6x7_subscript1_share1 , x2x4x5x6_subscript1_share1 , x2x4x5x7_subscript1_share1 , x2x4x6x7_subscript1_share1 , x2x5x6x7_subscript1_share1 , x3x4x5x6_subscript1_share1 , x3x4x5x7_subscript1_share1 , x3x4x6x7_subscript1_share1 , x3x5x6x7_subscript1_share1 , x4x5x6x7_subscript1_share1 , x0x1x2x3x4_subscript1_share1 , x0x1x2x3x5_subscript1_share1 , x0x1x2x3x6_subscript1_share1 , x0x1x2x3x7_subscript1_share1 , x0x1x2x4x5_subscript1_share1 , x0x1x2x4x6_subscript1_share1 , x0x1x2x4x7_subscript1_share1 , x0x1x2x5x6_subscript1_share1 , x0x1x2x5x7_subscript1_share1 , x0x1x2x6x7_subscript1_share1 , x0x1x3x4x5_subscript1_share1 , x0x1x3x4x6_subscript1_share1 , x0x1x3x4x7_subscript1_share1 , x0x1x3x5x6_subscript1_share1 , x0x1x3x5x7_subscript1_share1 , x0x1x3x6x7_subscript1_share1 , x0x1x4x5x6_subscript1_share1 , x0x1x4x5x7_subscript1_share1 , x0x1x4x6x7_subscript1_share1 , x0x1x5x6x7_subscript1_share1 , x0x2x3x4x5_subscript1_share1 , x0x2x3x4x6_subscript1_share1 , x0x2x3x4x7_subscript1_share1 , x0x2x3x5x6_subscript1_share1 , x0x2x3x5x7_subscript1_share1 , x0x2x3x6x7_subscript1_share1 , x0x2x4x5x6_subscript1_share1 , x0x2x4x5x7_subscript1_share1 , x0x2x4x6x7_subscript1_share1 , x0x2x5x6x7_subscript1_share1 , x0x3x4x5x6_subscript1_share1 , x0x3x4x5x7_subscript1_share1 , x0x3x4x6x7_subscript1_share1 , x0x3x5x6x7_subscript1_share1 , x0x4x5x6x7_subscript1_share1 , x1x2x3x4x5_subscript1_share1 , x1x2x3x4x6_subscript1_share1 , x1x2x3x4x7_subscript1_share1 , x1x2x3x5x6_subscript1_share1 , x1x2x3x5x7_subscript1_share1 , x1x2x3x6x7_subscript1_share1 , x1x2x4x5x6_subscript1_share1 , x1x2x4x5x7_subscript1_share1 , x1x2x4x6x7_subscript1_share1 , x1x2x5x6x7_subscript1_share1 , x1x3x4x5x6_subscript1_share1 , x1x3x4x5x7_subscript1_share1 , x1x3x4x6x7_subscript1_share1 , x1x3x5x6x7_subscript1_share1 , x1x4x5x6x7_subscript1_share1 , x2x3x4x5x6_subscript1_share1 , x2x3x4x5x7_subscript1_share1 , x2x3x4x6x7_subscript1_share1 , x2x3x5x6x7_subscript1_share1 , x2x4x5x6x7_subscript1_share1 , x3x4x5x6x7_subscript1_share1 , x0x1x2x3x4x5_subscript1_share1 , x0x1x2x3x4x6_subscript1_share1 , x0x1x2x3x4x7_subscript1_share1 , x0x1x2x3x5x6_subscript1_share1 , x0x1x2x3x5x7_subscript1_share1 , x0x1x2x3x6x7_subscript1_share1 , x0x1x2x4x5x6_subscript1_share1 , x0x1x2x4x5x7_subscript1_share1 , x0x1x2x4x6x7_subscript1_share1 , x0x1x2x5x6x7_subscript1_share1 , x0x1x3x4x5x6_subscript1_share1 , x0x1x3x4x5x7_subscript1_share1 , x0x1x3x4x6x7_subscript1_share1 , x0x1x3x5x6x7_subscript1_share1 , x0x1x4x5x6x7_subscript1_share1 , x0x2x3x4x5x6_subscript1_share1 , x0x2x3x4x5x7_subscript1_share1 , x0x2x3x4x6x7_subscript1_share1 , x0x2x3x5x6x7_subscript1_share1 , x0x2x4x5x6x7_subscript1_share1 , x0x3x4x5x6x7_subscript1_share1 , x1x2x3x4x5x6_subscript1_share1 , x1x2x3x4x5x7_subscript1_share1 , x1x2x3x4x6x7_subscript1_share1 , x1x2x3x5x6x7_subscript1_share1 , x1x2x4x5x6x7_subscript1_share1 , x1x3x4x5x6x7_subscript1_share1 , x2x3x4x5x6x7_subscript1_share1 , x0x1x2x3x4x5x6_subscript1_share1 , x0x1x2x3x4x5x7_subscript1_share1 , x0x1x2x3x4x6x7_subscript1_share1 , x0x1x2x3x5x6x7_subscript1_share1 , x0x1x2x4x5x6x7_subscript1_share1 , x0x1x3x4x5x6x7_subscript1_share1 , x0x2x3x4x5x6x7_subscript1_share1 , x1x2x3x4x5x6x7_subscript1_share1 
);

combi_logic_cycle2_output_share2 inst_second_cycle_share2(
    x0_subscript0_share2_reg , x2_subscript0_share2_reg , x3_subscript0_share2_reg , x4_subscript0_share2_reg , x6_subscript0_share2_reg , x7_subscript0_share2_reg , x1_subscript0_share2_reg , x5_subscript0_share2_reg , x0x1_subscript0_share2_reg , x0x4_subscript0_share2_reg , x0x5_subscript0_share2_reg , x0x6_subscript0_share2_reg , x1x2_subscript0_share2_reg , x1x3_subscript0_share2_reg , x1x4_subscript0_share2_reg , x1x6_subscript0_share2_reg , x2x3_subscript0_share2_reg , x2x4_subscript0_share2_reg , x2x6_subscript0_share2_reg , x2x7_subscript0_share2_reg , x4x6_subscript0_share2_reg , x5x6_subscript0_share2_reg , x5x7_subscript0_share2_reg , x6x7_subscript0_share2_reg , x0x2_subscript0_share2_reg , x0x3_subscript0_share2_reg , x0x7_subscript0_share2_reg , x1x7_subscript0_share2_reg , x3x7_subscript0_share2_reg , x4x5_subscript0_share2_reg , x3x4_subscript0_share2_reg , x4x7_subscript0_share2_reg , x3x6_subscript0_share2_reg , x1x5_subscript0_share2_reg , x2x5_subscript0_share2_reg , x3x5_subscript0_share2_reg , x0x1x4_subscript0_share2_reg , x0x1x6_subscript0_share2_reg , x0x1x7_subscript0_share2_reg , x0x2x4_subscript0_share2_reg , x0x2x5_subscript0_share2_reg , x0x2x6_subscript0_share2_reg , x0x2x7_subscript0_share2_reg , x0x3x4_subscript0_share2_reg , x0x3x5_subscript0_share2_reg , x0x3x6_subscript0_share2_reg , x0x4x6_subscript0_share2_reg , x0x4x7_subscript0_share2_reg , x1x2x3_subscript0_share2_reg , x1x2x4_subscript0_share2_reg , x1x2x6_subscript0_share2_reg , x1x3x4_subscript0_share2_reg , x1x3x7_subscript0_share2_reg , x1x4x6_subscript0_share2_reg , x1x5x6_subscript0_share2_reg , x2x3x5_subscript0_share2_reg , x2x3x7_subscript0_share2_reg , x2x4x7_subscript0_share2_reg , x2x5x6_subscript0_share2_reg , x2x5x7_subscript0_share2_reg , x2x6x7_subscript0_share2_reg , x3x4x7_subscript0_share2_reg , x3x5x7_subscript0_share2_reg , x3x6x7_subscript0_share2_reg , x4x5x6_subscript0_share2_reg , x5x6x7_subscript0_share2_reg , x0x1x3_subscript0_share2_reg , x0x2x3_subscript0_share2_reg , x0x4x5_subscript0_share2_reg , x0x5x7_subscript0_share2_reg , x0x6x7_subscript0_share2_reg , x1x3x5_subscript0_share2_reg , x1x3x6_subscript0_share2_reg , x1x4x7_subscript0_share2_reg , x2x3x4_subscript0_share2_reg , x2x3x6_subscript0_share2_reg , x3x4x6_subscript0_share2_reg , x3x5x6_subscript0_share2_reg , x0x1x5_subscript0_share2_reg , x0x3x7_subscript0_share2_reg , x1x2x5_subscript0_share2_reg , x1x2x7_subscript0_share2_reg , x1x4x5_subscript0_share2_reg , x1x5x7_subscript0_share2_reg , x2x4x5_subscript0_share2_reg , x3x4x5_subscript0_share2_reg , x4x6x7_subscript0_share2_reg , x1x6x7_subscript0_share2_reg , x4x5x7_subscript0_share2_reg , x0x1x2_subscript0_share2_reg , x0x5x6_subscript0_share2_reg , x2x4x6_subscript0_share2_reg , x0x1x2x3_subscript0_share2_reg , x0x1x2x5_subscript0_share2_reg , x0x1x2x6_subscript0_share2_reg , x0x1x2x7_subscript0_share2_reg , x0x1x4x5_subscript0_share2_reg , x0x1x4x7_subscript0_share2_reg , x0x2x3x5_subscript0_share2_reg , x0x2x3x7_subscript0_share2_reg , x0x2x4x5_subscript0_share2_reg , x0x2x4x7_subscript0_share2_reg , x0x2x5x6_subscript0_share2_reg , x0x2x5x7_subscript0_share2_reg , x0x3x4x6_subscript0_share2_reg , x0x3x5x6_subscript0_share2_reg , x0x4x5x6_subscript0_share2_reg , x0x4x5x7_subscript0_share2_reg , x0x4x6x7_subscript0_share2_reg , x1x2x3x5_subscript0_share2_reg , x1x2x3x6_subscript0_share2_reg , x1x2x3x7_subscript0_share2_reg , x1x2x4x6_subscript0_share2_reg , x1x2x4x7_subscript0_share2_reg , x1x2x6x7_subscript0_share2_reg , x1x3x4x6_subscript0_share2_reg , x1x3x6x7_subscript0_share2_reg , x1x4x5x6_subscript0_share2_reg , x1x4x5x7_subscript0_share2_reg , x1x5x6x7_subscript0_share2_reg , x2x3x5x7_subscript0_share2_reg , x2x3x6x7_subscript0_share2_reg , x2x4x5x6_subscript0_share2_reg , x2x4x5x7_subscript0_share2_reg , x3x5x6x7_subscript0_share2_reg , x0x1x3x4_subscript0_share2_reg , x0x1x3x6_subscript0_share2_reg , x0x1x5x6_subscript0_share2_reg , x0x2x3x6_subscript0_share2_reg , x0x3x4x5_subscript0_share2_reg , x1x2x5x6_subscript0_share2_reg , x1x2x5x7_subscript0_share2_reg , x1x3x4x5_subscript0_share2_reg , x1x3x4x7_subscript0_share2_reg , x1x3x5x6_subscript0_share2_reg , x1x3x5x7_subscript0_share2_reg , x1x4x6x7_subscript0_share2_reg , x2x3x4x5_subscript0_share2_reg , x2x3x4x7_subscript0_share2_reg , x2x4x6x7_subscript0_share2_reg , x3x4x5x6_subscript0_share2_reg , x3x4x5x7_subscript0_share2_reg , x3x4x6x7_subscript0_share2_reg , x0x1x3x5_subscript0_share2_reg , x0x1x4x6_subscript0_share2_reg , x0x2x3x4_subscript0_share2_reg , x0x2x4x6_subscript0_share2_reg , x0x3x4x7_subscript0_share2_reg , x0x3x5x7_subscript0_share2_reg , x1x2x3x4_subscript0_share2_reg , x2x3x4x6_subscript0_share2_reg , x2x3x5x6_subscript0_share2_reg , x2x5x6x7_subscript0_share2_reg , x4x5x6x7_subscript0_share2_reg , x0x1x2x4_subscript0_share2_reg , x0x1x6x7_subscript0_share2_reg , x0x2x6x7_subscript0_share2_reg , x0x3x6x7_subscript0_share2_reg , x0x5x6x7_subscript0_share2_reg , x1x2x4x5_subscript0_share2_reg , x0x1x3x7_subscript0_share2_reg , x0x1x5x7_subscript0_share2_reg , x0x1x2x3x4_subscript0_share2_reg , x0x1x2x3x6_subscript0_share2_reg , x0x1x2x3x7_subscript0_share2_reg , x0x1x2x4x5_subscript0_share2_reg , x0x1x2x4x7_subscript0_share2_reg , x0x1x2x5x7_subscript0_share2_reg , x0x1x2x6x7_subscript0_share2_reg , x0x1x3x4x6_subscript0_share2_reg , x0x1x3x5x6_subscript0_share2_reg , x0x1x3x5x7_subscript0_share2_reg , x0x1x3x6x7_subscript0_share2_reg , x0x1x4x5x6_subscript0_share2_reg , x0x1x5x6x7_subscript0_share2_reg , x0x2x3x4x5_subscript0_share2_reg , x0x2x3x4x6_subscript0_share2_reg , x0x2x4x5x7_subscript0_share2_reg , x0x2x4x6x7_subscript0_share2_reg , x0x3x4x5x6_subscript0_share2_reg , x0x3x4x5x7_subscript0_share2_reg , x0x3x4x6x7_subscript0_share2_reg , x0x3x5x6x7_subscript0_share2_reg , x1x2x3x5x6_subscript0_share2_reg , x1x2x3x5x7_subscript0_share2_reg , x1x2x4x5x6_subscript0_share2_reg , x1x2x4x6x7_subscript0_share2_reg , x1x2x5x6x7_subscript0_share2_reg , x1x3x4x5x7_subscript0_share2_reg , x2x3x4x5x6_subscript0_share2_reg , x2x3x4x5x7_subscript0_share2_reg , x2x4x5x6x7_subscript0_share2_reg , x0x1x2x4x6_subscript0_share2_reg , x0x1x3x4x7_subscript0_share2_reg , x0x2x3x4x7_subscript0_share2_reg , x0x2x3x5x7_subscript0_share2_reg , x0x2x3x6x7_subscript0_share2_reg , x0x2x4x5x6_subscript0_share2_reg , x0x2x5x6x7_subscript0_share2_reg , x0x4x5x6x7_subscript0_share2_reg , x1x2x3x4x6_subscript0_share2_reg , x1x3x4x5x6_subscript0_share2_reg , x2x3x4x6x7_subscript0_share2_reg , x0x1x2x3x5_subscript0_share2_reg , x0x1x4x6x7_subscript0_share2_reg , x1x2x3x4x5_subscript0_share2_reg , x1x2x3x6x7_subscript0_share2_reg , x1x2x4x5x7_subscript0_share2_reg , x1x3x4x6x7_subscript0_share2_reg , x1x3x5x6x7_subscript0_share2_reg , x1x4x5x6x7_subscript0_share2_reg , x2x3x5x6x7_subscript0_share2_reg , x3x4x5x6x7_subscript0_share2_reg , x0x1x2x5x6_subscript0_share2_reg , x0x1x3x4x5_subscript0_share2_reg , x0x1x4x5x7_subscript0_share2_reg , x0x2x3x5x6_subscript0_share2_reg , x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x4x6_subscript0_share2_reg , x0x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x5x7_subscript0_share2_reg , x0x1x2x3x6x7_subscript0_share2_reg , x0x1x2x4x5x7_subscript0_share2_reg , x0x1x2x5x6x7_subscript0_share2_reg , x0x1x3x4x6x7_subscript0_share2_reg , x0x1x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6_subscript0_share2_reg , x0x2x3x4x5x7_subscript0_share2_reg , x0x2x3x5x6x7_subscript0_share2_reg , x1x2x3x4x6x7_subscript0_share2_reg , x1x2x4x5x6x7_subscript0_share2_reg , x1x3x4x5x6x7_subscript0_share2_reg , x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6_subscript0_share2_reg , x0x1x2x4x6x7_subscript0_share2_reg , x0x1x3x4x5x6_subscript0_share2_reg , x0x2x3x4x6x7_subscript0_share2_reg , x1x2x3x4x5x6_subscript0_share2_reg , x1x2x3x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5_subscript0_share2_reg , x0x1x2x4x5x6_subscript0_share2_reg , x0x1x3x4x5x7_subscript0_share2_reg , x0x1x3x5x6x7_subscript0_share2_reg , x0x2x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x7_subscript0_share2_reg , x0x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x6x7_subscript0_share2_reg , x0x1x2x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6x7_subscript0_share2_reg , x0x1x3x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5x6_subscript0_share2_reg , x0x1x2x3x4x5x7_subscript0_share2_reg , 
    x0_pipelined_share2_reg ,x1_pipelined_share2_reg ,x2_pipelined_share2_reg ,x3_pipelined_share2_reg ,x4_pipelined_share2_reg ,x5_pipelined_share2_reg ,x6_pipelined_share2_reg ,x7_pipelined_share2_reg ,
    x0_subscript1_share2, x1_subscript1_share2, x2_subscript1_share2, x3_subscript1_share2, x4_subscript1_share2, x5_subscript1_share2, x6_subscript1_share2, x7_subscript1_share2 , x0x1_subscript1_share2 , x0x2_subscript1_share2 , x0x3_subscript1_share2 , x0x4_subscript1_share2 , x0x5_subscript1_share2 , x0x6_subscript1_share2 , x0x7_subscript1_share2 , x1x2_subscript1_share2 , x1x3_subscript1_share2 , x1x4_subscript1_share2 , x1x5_subscript1_share2 , x1x6_subscript1_share2 , x1x7_subscript1_share2 , x2x3_subscript1_share2 , x2x4_subscript1_share2 , x2x5_subscript1_share2 , x2x6_subscript1_share2 , x2x7_subscript1_share2 , x3x4_subscript1_share2 , x3x5_subscript1_share2 , x3x6_subscript1_share2 , x3x7_subscript1_share2 , x4x5_subscript1_share2 , x4x6_subscript1_share2 , x4x7_subscript1_share2 , x5x6_subscript1_share2 , x5x7_subscript1_share2 , x6x7_subscript1_share2 , x0x1x2_subscript1_share2 , x0x1x3_subscript1_share2 , x0x1x4_subscript1_share2 , x0x1x5_subscript1_share2 , x0x1x6_subscript1_share2 , x0x1x7_subscript1_share2 , x0x2x3_subscript1_share2 , x0x2x4_subscript1_share2 , x0x2x5_subscript1_share2 , x0x2x6_subscript1_share2 , x0x2x7_subscript1_share2 , x0x3x4_subscript1_share2 , x0x3x5_subscript1_share2 , x0x3x6_subscript1_share2 , x0x3x7_subscript1_share2 , x0x4x5_subscript1_share2 , x0x4x6_subscript1_share2 , x0x4x7_subscript1_share2 , x0x5x6_subscript1_share2 , x0x5x7_subscript1_share2 , x0x6x7_subscript1_share2 , x1x2x3_subscript1_share2 , x1x2x4_subscript1_share2 , x1x2x5_subscript1_share2 , x1x2x6_subscript1_share2 , x1x2x7_subscript1_share2 , x1x3x4_subscript1_share2 , x1x3x5_subscript1_share2 , x1x3x6_subscript1_share2 , x1x3x7_subscript1_share2 , x1x4x5_subscript1_share2 , x1x4x6_subscript1_share2 , x1x4x7_subscript1_share2 , x1x5x6_subscript1_share2 , x1x5x7_subscript1_share2 , x1x6x7_subscript1_share2 , x2x3x4_subscript1_share2 , x2x3x5_subscript1_share2 , x2x3x6_subscript1_share2 , x2x3x7_subscript1_share2 , x2x4x5_subscript1_share2 , x2x4x6_subscript1_share2 , x2x4x7_subscript1_share2 , x2x5x6_subscript1_share2 , x2x5x7_subscript1_share2 , x2x6x7_subscript1_share2 , x3x4x5_subscript1_share2 , x3x4x6_subscript1_share2 , x3x4x7_subscript1_share2 , x3x5x6_subscript1_share2 , x3x5x7_subscript1_share2 , x3x6x7_subscript1_share2 , x4x5x6_subscript1_share2 , x4x5x7_subscript1_share2 , x4x6x7_subscript1_share2 , x5x6x7_subscript1_share2 , x0x1x2x3_subscript1_share2 , x0x1x2x4_subscript1_share2 , x0x1x2x5_subscript1_share2 , x0x1x2x6_subscript1_share2 , x0x1x2x7_subscript1_share2 , x0x1x3x4_subscript1_share2 , x0x1x3x5_subscript1_share2 , x0x1x3x6_subscript1_share2 , x0x1x3x7_subscript1_share2 , x0x1x4x5_subscript1_share2 , x0x1x4x6_subscript1_share2 , x0x1x4x7_subscript1_share2 , x0x1x5x6_subscript1_share2 , x0x1x5x7_subscript1_share2 , x0x1x6x7_subscript1_share2 , x0x2x3x4_subscript1_share2 , x0x2x3x5_subscript1_share2 , x0x2x3x6_subscript1_share2 , x0x2x3x7_subscript1_share2 , x0x2x4x5_subscript1_share2 , x0x2x4x6_subscript1_share2 , x0x2x4x7_subscript1_share2 , x0x2x5x6_subscript1_share2 , x0x2x5x7_subscript1_share2 , x0x2x6x7_subscript1_share2 , x0x3x4x5_subscript1_share2 , x0x3x4x6_subscript1_share2 , x0x3x4x7_subscript1_share2 , x0x3x5x6_subscript1_share2 , x0x3x5x7_subscript1_share2 , x0x3x6x7_subscript1_share2 , x0x4x5x6_subscript1_share2 , x0x4x5x7_subscript1_share2 , x0x4x6x7_subscript1_share2 , x0x5x6x7_subscript1_share2 , x1x2x3x4_subscript1_share2 , x1x2x3x5_subscript1_share2 , x1x2x3x6_subscript1_share2 , x1x2x3x7_subscript1_share2 , x1x2x4x5_subscript1_share2 , x1x2x4x6_subscript1_share2 , x1x2x4x7_subscript1_share2 , x1x2x5x6_subscript1_share2 , x1x2x5x7_subscript1_share2 , x1x2x6x7_subscript1_share2 , x1x3x4x5_subscript1_share2 , x1x3x4x6_subscript1_share2 , x1x3x4x7_subscript1_share2 , x1x3x5x6_subscript1_share2 , x1x3x5x7_subscript1_share2 , x1x3x6x7_subscript1_share2 , x1x4x5x6_subscript1_share2 , x1x4x5x7_subscript1_share2 , x1x4x6x7_subscript1_share2 , x1x5x6x7_subscript1_share2 , x2x3x4x5_subscript1_share2 , x2x3x4x6_subscript1_share2 , x2x3x4x7_subscript1_share2 , x2x3x5x6_subscript1_share2 , x2x3x5x7_subscript1_share2 , x2x3x6x7_subscript1_share2 , x2x4x5x6_subscript1_share2 , x2x4x5x7_subscript1_share2 , x2x4x6x7_subscript1_share2 , x2x5x6x7_subscript1_share2 , x3x4x5x6_subscript1_share2 , x3x4x5x7_subscript1_share2 , x3x4x6x7_subscript1_share2 , x3x5x6x7_subscript1_share2 , x4x5x6x7_subscript1_share2 , x0x1x2x3x4_subscript1_share2 , x0x1x2x3x5_subscript1_share2 , x0x1x2x3x6_subscript1_share2 , x0x1x2x3x7_subscript1_share2 , x0x1x2x4x5_subscript1_share2 , x0x1x2x4x6_subscript1_share2 , x0x1x2x4x7_subscript1_share2 , x0x1x2x5x6_subscript1_share2 , x0x1x2x5x7_subscript1_share2 , x0x1x2x6x7_subscript1_share2 , x0x1x3x4x5_subscript1_share2 , x0x1x3x4x6_subscript1_share2 , x0x1x3x4x7_subscript1_share2 , x0x1x3x5x6_subscript1_share2 , x0x1x3x5x7_subscript1_share2 , x0x1x3x6x7_subscript1_share2 , x0x1x4x5x6_subscript1_share2 , x0x1x4x5x7_subscript1_share2 , x0x1x4x6x7_subscript1_share2 , x0x1x5x6x7_subscript1_share2 , x0x2x3x4x5_subscript1_share2 , x0x2x3x4x6_subscript1_share2 , x0x2x3x4x7_subscript1_share2 , x0x2x3x5x6_subscript1_share2 , x0x2x3x5x7_subscript1_share2 , x0x2x3x6x7_subscript1_share2 , x0x2x4x5x6_subscript1_share2 , x0x2x4x5x7_subscript1_share2 , x0x2x4x6x7_subscript1_share2 , x0x2x5x6x7_subscript1_share2 , x0x3x4x5x6_subscript1_share2 , x0x3x4x5x7_subscript1_share2 , x0x3x4x6x7_subscript1_share2 , x0x3x5x6x7_subscript1_share2 , x0x4x5x6x7_subscript1_share2 , x1x2x3x4x5_subscript1_share2 , x1x2x3x4x6_subscript1_share2 , x1x2x3x4x7_subscript1_share2 , x1x2x3x5x6_subscript1_share2 , x1x2x3x5x7_subscript1_share2 , x1x2x3x6x7_subscript1_share2 , x1x2x4x5x6_subscript1_share2 , x1x2x4x5x7_subscript1_share2 , x1x2x4x6x7_subscript1_share2 , x1x2x5x6x7_subscript1_share2 , x1x3x4x5x6_subscript1_share2 , x1x3x4x5x7_subscript1_share2 , x1x3x4x6x7_subscript1_share2 , x1x3x5x6x7_subscript1_share2 , x1x4x5x6x7_subscript1_share2 , x2x3x4x5x6_subscript1_share2 , x2x3x4x5x7_subscript1_share2 , x2x3x4x6x7_subscript1_share2 , x2x3x5x6x7_subscript1_share2 , x2x4x5x6x7_subscript1_share2 , x3x4x5x6x7_subscript1_share2 , x0x1x2x3x4x5_subscript1_share2 , x0x1x2x3x4x6_subscript1_share2 , x0x1x2x3x4x7_subscript1_share2 , x0x1x2x3x5x6_subscript1_share2 , x0x1x2x3x5x7_subscript1_share2 , x0x1x2x3x6x7_subscript1_share2 , x0x1x2x4x5x6_subscript1_share2 , x0x1x2x4x5x7_subscript1_share2 , x0x1x2x4x6x7_subscript1_share2 , x0x1x2x5x6x7_subscript1_share2 , x0x1x3x4x5x6_subscript1_share2 , x0x1x3x4x5x7_subscript1_share2 , x0x1x3x4x6x7_subscript1_share2 , x0x1x3x5x6x7_subscript1_share2 , x0x1x4x5x6x7_subscript1_share2 , x0x2x3x4x5x6_subscript1_share2 , x0x2x3x4x5x7_subscript1_share2 , x0x2x3x4x6x7_subscript1_share2 , x0x2x3x5x6x7_subscript1_share2 , x0x2x4x5x6x7_subscript1_share2 , x0x3x4x5x6x7_subscript1_share2 , x1x2x3x4x5x6_subscript1_share2 , x1x2x3x4x5x7_subscript1_share2 , x1x2x3x4x6x7_subscript1_share2 , x1x2x3x5x6x7_subscript1_share2 , x1x2x4x5x6x7_subscript1_share2 , x1x3x4x5x6x7_subscript1_share2 , x2x3x4x5x6x7_subscript1_share2 , x0x1x2x3x4x5x6_subscript1_share2 , x0x1x2x3x4x5x7_subscript1_share2 , x0x1x2x3x4x6x7_subscript1_share2 , x0x1x2x3x5x6x7_subscript1_share2 , x0x1x2x4x5x6x7_subscript1_share2 , x0x1x3x4x5x6x7_subscript1_share2 , x0x2x3x4x5x6x7_subscript1_share2 , x1x2x3x4x5x6x7_subscript1_share2 
);


wire [254:1] rand_second_cycle_a ;
assign rand_second_cycle_a = rand_bit_cycle2[254:1];
wire [254:1] rand_second_cycle_b ;
assign rand_second_cycle_b = rand_bit_cycle2[508:255];

xor_AES_twofiftyfour xor_second_cycle_first_share(
    x0_subscript1_share1, x1_subscript1_share1, x2_subscript1_share1, x3_subscript1_share1, x4_subscript1_share1, x5_subscript1_share1, x6_subscript1_share1, x7_subscript1_share1 , x0x1_subscript1_share1 , x0x2_subscript1_share1 , x0x3_subscript1_share1 , x0x4_subscript1_share1 , x0x5_subscript1_share1 , x0x6_subscript1_share1 , x0x7_subscript1_share1 , x1x2_subscript1_share1 , x1x3_subscript1_share1 , x1x4_subscript1_share1 , x1x5_subscript1_share1 , x1x6_subscript1_share1 , x1x7_subscript1_share1 , x2x3_subscript1_share1 , x2x4_subscript1_share1 , x2x5_subscript1_share1 , x2x6_subscript1_share1 , x2x7_subscript1_share1 , x3x4_subscript1_share1 , x3x5_subscript1_share1 , x3x6_subscript1_share1 , x3x7_subscript1_share1 , x4x5_subscript1_share1 , x4x6_subscript1_share1 , x4x7_subscript1_share1 , x5x6_subscript1_share1 , x5x7_subscript1_share1 , x6x7_subscript1_share1 , x0x1x2_subscript1_share1 , x0x1x3_subscript1_share1 , x0x1x4_subscript1_share1 , x0x1x5_subscript1_share1 , x0x1x6_subscript1_share1 , x0x1x7_subscript1_share1 , x0x2x3_subscript1_share1 , x0x2x4_subscript1_share1 , x0x2x5_subscript1_share1 , x0x2x6_subscript1_share1 , x0x2x7_subscript1_share1 , x0x3x4_subscript1_share1 , x0x3x5_subscript1_share1 , x0x3x6_subscript1_share1 , x0x3x7_subscript1_share1 , x0x4x5_subscript1_share1 , x0x4x6_subscript1_share1 , x0x4x7_subscript1_share1 , x0x5x6_subscript1_share1 , x0x5x7_subscript1_share1 , x0x6x7_subscript1_share1 , x1x2x3_subscript1_share1 , x1x2x4_subscript1_share1 , x1x2x5_subscript1_share1 , x1x2x6_subscript1_share1 , x1x2x7_subscript1_share1 , x1x3x4_subscript1_share1 , x1x3x5_subscript1_share1 , x1x3x6_subscript1_share1 , x1x3x7_subscript1_share1 , x1x4x5_subscript1_share1 , x1x4x6_subscript1_share1 , x1x4x7_subscript1_share1 , x1x5x6_subscript1_share1 , x1x5x7_subscript1_share1 , x1x6x7_subscript1_share1 , x2x3x4_subscript1_share1 , x2x3x5_subscript1_share1 , x2x3x6_subscript1_share1 , x2x3x7_subscript1_share1 , x2x4x5_subscript1_share1 , x2x4x6_subscript1_share1 , x2x4x7_subscript1_share1 , x2x5x6_subscript1_share1 , x2x5x7_subscript1_share1 , x2x6x7_subscript1_share1 , x3x4x5_subscript1_share1 , x3x4x6_subscript1_share1 , x3x4x7_subscript1_share1 , x3x5x6_subscript1_share1 , x3x5x7_subscript1_share1 , x3x6x7_subscript1_share1 , x4x5x6_subscript1_share1 , x4x5x7_subscript1_share1 , x4x6x7_subscript1_share1 , x5x6x7_subscript1_share1 , x0x1x2x3_subscript1_share1 , x0x1x2x4_subscript1_share1 , x0x1x2x5_subscript1_share1 , x0x1x2x6_subscript1_share1 , x0x1x2x7_subscript1_share1 , x0x1x3x4_subscript1_share1 , x0x1x3x5_subscript1_share1 , x0x1x3x6_subscript1_share1 , x0x1x3x7_subscript1_share1 , x0x1x4x5_subscript1_share1 , x0x1x4x6_subscript1_share1 , x0x1x4x7_subscript1_share1 , x0x1x5x6_subscript1_share1 , x0x1x5x7_subscript1_share1 , x0x1x6x7_subscript1_share1 , x0x2x3x4_subscript1_share1 , x0x2x3x5_subscript1_share1 , x0x2x3x6_subscript1_share1 , x0x2x3x7_subscript1_share1 , x0x2x4x5_subscript1_share1 , x0x2x4x6_subscript1_share1 , x0x2x4x7_subscript1_share1 , x0x2x5x6_subscript1_share1 , x0x2x5x7_subscript1_share1 , x0x2x6x7_subscript1_share1 , x0x3x4x5_subscript1_share1 , x0x3x4x6_subscript1_share1 , x0x3x4x7_subscript1_share1 , x0x3x5x6_subscript1_share1 , x0x3x5x7_subscript1_share1 , x0x3x6x7_subscript1_share1 , x0x4x5x6_subscript1_share1 , x0x4x5x7_subscript1_share1 , x0x4x6x7_subscript1_share1 , x0x5x6x7_subscript1_share1 , x1x2x3x4_subscript1_share1 , x1x2x3x5_subscript1_share1 , x1x2x3x6_subscript1_share1 , x1x2x3x7_subscript1_share1 , x1x2x4x5_subscript1_share1 , x1x2x4x6_subscript1_share1 , x1x2x4x7_subscript1_share1 , x1x2x5x6_subscript1_share1 , x1x2x5x7_subscript1_share1 , x1x2x6x7_subscript1_share1 , x1x3x4x5_subscript1_share1 , x1x3x4x6_subscript1_share1 , x1x3x4x7_subscript1_share1 , x1x3x5x6_subscript1_share1 , x1x3x5x7_subscript1_share1 , x1x3x6x7_subscript1_share1 , x1x4x5x6_subscript1_share1 , x1x4x5x7_subscript1_share1 , x1x4x6x7_subscript1_share1 , x1x5x6x7_subscript1_share1 , x2x3x4x5_subscript1_share1 , x2x3x4x6_subscript1_share1 , x2x3x4x7_subscript1_share1 , x2x3x5x6_subscript1_share1 , x2x3x5x7_subscript1_share1 , x2x3x6x7_subscript1_share1 , x2x4x5x6_subscript1_share1 , x2x4x5x7_subscript1_share1 , x2x4x6x7_subscript1_share1 , x2x5x6x7_subscript1_share1 , x3x4x5x6_subscript1_share1 , x3x4x5x7_subscript1_share1 , x3x4x6x7_subscript1_share1 , x3x5x6x7_subscript1_share1 , x4x5x6x7_subscript1_share1 , x0x1x2x3x4_subscript1_share1 , x0x1x2x3x5_subscript1_share1 , x0x1x2x3x6_subscript1_share1 , x0x1x2x3x7_subscript1_share1 , x0x1x2x4x5_subscript1_share1 , x0x1x2x4x6_subscript1_share1 , x0x1x2x4x7_subscript1_share1 , x0x1x2x5x6_subscript1_share1 , x0x1x2x5x7_subscript1_share1 , x0x1x2x6x7_subscript1_share1 , x0x1x3x4x5_subscript1_share1 , x0x1x3x4x6_subscript1_share1 , x0x1x3x4x7_subscript1_share1 , x0x1x3x5x6_subscript1_share1 , x0x1x3x5x7_subscript1_share1 , x0x1x3x6x7_subscript1_share1 , x0x1x4x5x6_subscript1_share1 , x0x1x4x5x7_subscript1_share1 , x0x1x4x6x7_subscript1_share1 , x0x1x5x6x7_subscript1_share1 , x0x2x3x4x5_subscript1_share1 , x0x2x3x4x6_subscript1_share1 , x0x2x3x4x7_subscript1_share1 , x0x2x3x5x6_subscript1_share1 , x0x2x3x5x7_subscript1_share1 , x0x2x3x6x7_subscript1_share1 , x0x2x4x5x6_subscript1_share1 , x0x2x4x5x7_subscript1_share1 , x0x2x4x6x7_subscript1_share1 , x0x2x5x6x7_subscript1_share1 , x0x3x4x5x6_subscript1_share1 , x0x3x4x5x7_subscript1_share1 , x0x3x4x6x7_subscript1_share1 , x0x3x5x6x7_subscript1_share1 , x0x4x5x6x7_subscript1_share1 , x1x2x3x4x5_subscript1_share1 , x1x2x3x4x6_subscript1_share1 , x1x2x3x4x7_subscript1_share1 , x1x2x3x5x6_subscript1_share1 , x1x2x3x5x7_subscript1_share1 , x1x2x3x6x7_subscript1_share1 , x1x2x4x5x6_subscript1_share1 , x1x2x4x5x7_subscript1_share1 , x1x2x4x6x7_subscript1_share1 , x1x2x5x6x7_subscript1_share1 , x1x3x4x5x6_subscript1_share1 , x1x3x4x5x7_subscript1_share1 , x1x3x4x6x7_subscript1_share1 , x1x3x5x6x7_subscript1_share1 , x1x4x5x6x7_subscript1_share1 , x2x3x4x5x6_subscript1_share1 , x2x3x4x5x7_subscript1_share1 , x2x3x4x6x7_subscript1_share1 , x2x3x5x6x7_subscript1_share1 , x2x4x5x6x7_subscript1_share1 , x3x4x5x6x7_subscript1_share1 , x0x1x2x3x4x5_subscript1_share1 , x0x1x2x3x4x6_subscript1_share1 , x0x1x2x3x4x7_subscript1_share1 , x0x1x2x3x5x6_subscript1_share1 , x0x1x2x3x5x7_subscript1_share1 , x0x1x2x3x6x7_subscript1_share1 , x0x1x2x4x5x6_subscript1_share1 , x0x1x2x4x5x7_subscript1_share1 , x0x1x2x4x6x7_subscript1_share1 , x0x1x2x5x6x7_subscript1_share1 , x0x1x3x4x5x6_subscript1_share1 , x0x1x3x4x5x7_subscript1_share1 , x0x1x3x4x6x7_subscript1_share1 , x0x1x3x5x6x7_subscript1_share1 , x0x1x4x5x6x7_subscript1_share1 , x0x2x3x4x5x6_subscript1_share1 , x0x2x3x4x5x7_subscript1_share1 , x0x2x3x4x6x7_subscript1_share1 , x0x2x3x5x6x7_subscript1_share1 , x0x2x4x5x6x7_subscript1_share1 , x0x3x4x5x6x7_subscript1_share1 , x1x2x3x4x5x6_subscript1_share1 , x1x2x3x4x5x7_subscript1_share1 , x1x2x3x4x6x7_subscript1_share1 , x1x2x3x5x6x7_subscript1_share1 , x1x2x4x5x6x7_subscript1_share1 , x1x3x4x5x6x7_subscript1_share1 , x2x3x4x5x6x7_subscript1_share1 , x0x1x2x3x4x5x6_subscript1_share1 , x0x1x2x3x4x5x7_subscript1_share1 , x0x1x2x3x4x6x7_subscript1_share1 , x0x1x2x3x5x6x7_subscript1_share1 , x0x1x2x4x5x6x7_subscript1_share1 , x0x1x3x4x5x6x7_subscript1_share1 , x0x2x3x4x5x6x7_subscript1_share1 , x1x2x3x4x5x6x7_subscript1_share1 ,
    rand_second_cycle_a[1] ,rand_second_cycle_a[2] ,rand_second_cycle_a[3] ,rand_second_cycle_a[4] ,rand_second_cycle_a[5] ,rand_second_cycle_a[6] ,rand_second_cycle_a[7] ,rand_second_cycle_a[8] ,rand_second_cycle_a[9] ,rand_second_cycle_a[10] ,rand_second_cycle_a[11] ,rand_second_cycle_a[12] ,rand_second_cycle_a[13] ,rand_second_cycle_a[14] ,rand_second_cycle_a[15] ,rand_second_cycle_a[16] ,rand_second_cycle_a[17] ,rand_second_cycle_a[18] ,rand_second_cycle_a[19] ,rand_second_cycle_a[20] ,rand_second_cycle_a[21] ,rand_second_cycle_a[22] ,rand_second_cycle_a[23] ,rand_second_cycle_a[24] ,rand_second_cycle_a[25] ,rand_second_cycle_a[26] ,rand_second_cycle_a[27] ,rand_second_cycle_a[28] ,rand_second_cycle_a[29] ,rand_second_cycle_a[30] ,rand_second_cycle_a[31] ,rand_second_cycle_a[32] ,rand_second_cycle_a[33] ,rand_second_cycle_a[34] ,rand_second_cycle_a[35] ,rand_second_cycle_a[36] ,rand_second_cycle_a[37] ,rand_second_cycle_a[38] ,rand_second_cycle_a[39] ,rand_second_cycle_a[40] ,rand_second_cycle_a[41] ,rand_second_cycle_a[42] ,rand_second_cycle_a[43] ,rand_second_cycle_a[44] ,rand_second_cycle_a[45] ,rand_second_cycle_a[46] ,rand_second_cycle_a[47] ,rand_second_cycle_a[48] ,rand_second_cycle_a[49] ,rand_second_cycle_a[50] ,rand_second_cycle_a[51] ,rand_second_cycle_a[52] ,rand_second_cycle_a[53] ,rand_second_cycle_a[54] ,rand_second_cycle_a[55] ,rand_second_cycle_a[56] ,rand_second_cycle_a[57] ,rand_second_cycle_a[58] ,rand_second_cycle_a[59] ,rand_second_cycle_a[60] ,rand_second_cycle_a[61] ,rand_second_cycle_a[62] ,rand_second_cycle_a[63] ,rand_second_cycle_a[64] ,rand_second_cycle_a[65] ,rand_second_cycle_a[66] ,rand_second_cycle_a[67] ,rand_second_cycle_a[68] ,rand_second_cycle_a[69] ,rand_second_cycle_a[70] ,rand_second_cycle_a[71] ,rand_second_cycle_a[72] ,rand_second_cycle_a[73] ,rand_second_cycle_a[74] ,rand_second_cycle_a[75] ,rand_second_cycle_a[76] ,rand_second_cycle_a[77] ,rand_second_cycle_a[78] ,rand_second_cycle_a[79] ,rand_second_cycle_a[80] ,rand_second_cycle_a[81] ,rand_second_cycle_a[82] ,rand_second_cycle_a[83] ,rand_second_cycle_a[84] ,rand_second_cycle_a[85] ,rand_second_cycle_a[86] ,rand_second_cycle_a[87] ,rand_second_cycle_a[88] ,rand_second_cycle_a[89] ,rand_second_cycle_a[90] ,rand_second_cycle_a[91] ,rand_second_cycle_a[92] ,rand_second_cycle_a[93] ,rand_second_cycle_a[94] ,rand_second_cycle_a[95] ,rand_second_cycle_a[96] ,rand_second_cycle_a[97] ,rand_second_cycle_a[98] ,rand_second_cycle_a[99] ,rand_second_cycle_a[100] ,rand_second_cycle_a[101] ,rand_second_cycle_a[102] ,rand_second_cycle_a[103] ,rand_second_cycle_a[104] ,rand_second_cycle_a[105] ,rand_second_cycle_a[106] ,rand_second_cycle_a[107] ,rand_second_cycle_a[108] ,rand_second_cycle_a[109] ,rand_second_cycle_a[110] ,rand_second_cycle_a[111] ,rand_second_cycle_a[112] ,rand_second_cycle_a[113] ,rand_second_cycle_a[114] ,rand_second_cycle_a[115] ,rand_second_cycle_a[116] ,rand_second_cycle_a[117] ,rand_second_cycle_a[118] ,rand_second_cycle_a[119] ,rand_second_cycle_a[120] ,rand_second_cycle_a[121] ,rand_second_cycle_a[122] ,rand_second_cycle_a[123] ,rand_second_cycle_a[124] ,rand_second_cycle_a[125] ,rand_second_cycle_a[126] ,rand_second_cycle_a[127] ,rand_second_cycle_a[128] ,rand_second_cycle_a[129] ,rand_second_cycle_a[130] ,rand_second_cycle_a[131] ,rand_second_cycle_a[132] ,rand_second_cycle_a[133] ,rand_second_cycle_a[134] ,rand_second_cycle_a[135] ,rand_second_cycle_a[136] ,rand_second_cycle_a[137] ,rand_second_cycle_a[138] ,rand_second_cycle_a[139] ,rand_second_cycle_a[140] ,rand_second_cycle_a[141] ,rand_second_cycle_a[142] ,rand_second_cycle_a[143] ,rand_second_cycle_a[144] ,rand_second_cycle_a[145] ,rand_second_cycle_a[146] ,rand_second_cycle_a[147] ,rand_second_cycle_a[148] ,rand_second_cycle_a[149] ,rand_second_cycle_a[150] ,rand_second_cycle_a[151] ,rand_second_cycle_a[152] ,rand_second_cycle_a[153] ,rand_second_cycle_a[154] ,rand_second_cycle_a[155] ,rand_second_cycle_a[156] ,rand_second_cycle_a[157] ,rand_second_cycle_a[158] ,rand_second_cycle_a[159] ,rand_second_cycle_a[160] ,rand_second_cycle_a[161] ,rand_second_cycle_a[162] ,rand_second_cycle_a[163] ,rand_second_cycle_a[164] ,rand_second_cycle_a[165] ,rand_second_cycle_a[166] ,rand_second_cycle_a[167] ,rand_second_cycle_a[168] ,rand_second_cycle_a[169] ,rand_second_cycle_a[170] ,rand_second_cycle_a[171] ,rand_second_cycle_a[172] ,rand_second_cycle_a[173] ,rand_second_cycle_a[174] ,rand_second_cycle_a[175] ,rand_second_cycle_a[176] ,rand_second_cycle_a[177] ,rand_second_cycle_a[178] ,rand_second_cycle_a[179] ,rand_second_cycle_a[180] ,rand_second_cycle_a[181] ,rand_second_cycle_a[182] ,rand_second_cycle_a[183] ,rand_second_cycle_a[184] ,rand_second_cycle_a[185] ,rand_second_cycle_a[186] ,rand_second_cycle_a[187] ,rand_second_cycle_a[188] ,rand_second_cycle_a[189] ,rand_second_cycle_a[190] ,rand_second_cycle_a[191] ,rand_second_cycle_a[192] ,rand_second_cycle_a[193] ,rand_second_cycle_a[194] ,rand_second_cycle_a[195] ,rand_second_cycle_a[196] ,rand_second_cycle_a[197] ,rand_second_cycle_a[198] ,rand_second_cycle_a[199] ,rand_second_cycle_a[200] ,rand_second_cycle_a[201] ,rand_second_cycle_a[202] ,rand_second_cycle_a[203] ,rand_second_cycle_a[204] ,rand_second_cycle_a[205] ,rand_second_cycle_a[206] ,rand_second_cycle_a[207] ,rand_second_cycle_a[208] ,rand_second_cycle_a[209] ,rand_second_cycle_a[210] ,rand_second_cycle_a[211] ,rand_second_cycle_a[212] ,rand_second_cycle_a[213] ,rand_second_cycle_a[214] ,rand_second_cycle_a[215] ,rand_second_cycle_a[216] ,rand_second_cycle_a[217] ,rand_second_cycle_a[218] ,rand_second_cycle_a[219] ,rand_second_cycle_a[220] ,rand_second_cycle_a[221] ,rand_second_cycle_a[222] ,rand_second_cycle_a[223] ,rand_second_cycle_a[224] ,rand_second_cycle_a[225] ,rand_second_cycle_a[226] ,rand_second_cycle_a[227] ,rand_second_cycle_a[228] ,rand_second_cycle_a[229] ,rand_second_cycle_a[230] ,rand_second_cycle_a[231] ,rand_second_cycle_a[232] ,rand_second_cycle_a[233] ,rand_second_cycle_a[234] ,rand_second_cycle_a[235] ,rand_second_cycle_a[236] ,rand_second_cycle_a[237] ,rand_second_cycle_a[238] ,rand_second_cycle_a[239] ,rand_second_cycle_a[240] ,rand_second_cycle_a[241] ,rand_second_cycle_a[242] ,rand_second_cycle_a[243] ,rand_second_cycle_a[244] ,rand_second_cycle_a[245] ,rand_second_cycle_a[246] ,rand_second_cycle_a[247] ,rand_second_cycle_a[248] ,rand_second_cycle_a[249] ,rand_second_cycle_a[250] ,rand_second_cycle_a[251] ,rand_second_cycle_a[252] ,rand_second_cycle_a[253] ,rand_second_cycle_a[254] ,
    x0_subscript1_share1_wire, x1_subscript1_share1_wire, x2_subscript1_share1_wire, x3_subscript1_share1_wire, x4_subscript1_share1_wire, x5_subscript1_share1_wire, x6_subscript1_share1_wire, x7_subscript1_share1_wire , x0x1_subscript1_share1_wire , x0x2_subscript1_share1_wire , x0x3_subscript1_share1_wire , x0x4_subscript1_share1_wire , x0x5_subscript1_share1_wire , x0x6_subscript1_share1_wire , x0x7_subscript1_share1_wire , x1x2_subscript1_share1_wire , x1x3_subscript1_share1_wire , x1x4_subscript1_share1_wire , x1x5_subscript1_share1_wire , x1x6_subscript1_share1_wire , x1x7_subscript1_share1_wire , x2x3_subscript1_share1_wire , x2x4_subscript1_share1_wire , x2x5_subscript1_share1_wire , x2x6_subscript1_share1_wire , x2x7_subscript1_share1_wire , x3x4_subscript1_share1_wire , x3x5_subscript1_share1_wire , x3x6_subscript1_share1_wire , x3x7_subscript1_share1_wire , x4x5_subscript1_share1_wire , x4x6_subscript1_share1_wire , x4x7_subscript1_share1_wire , x5x6_subscript1_share1_wire , x5x7_subscript1_share1_wire , x6x7_subscript1_share1_wire , x0x1x2_subscript1_share1_wire , x0x1x3_subscript1_share1_wire , x0x1x4_subscript1_share1_wire , x0x1x5_subscript1_share1_wire , x0x1x6_subscript1_share1_wire , x0x1x7_subscript1_share1_wire , x0x2x3_subscript1_share1_wire , x0x2x4_subscript1_share1_wire , x0x2x5_subscript1_share1_wire , x0x2x6_subscript1_share1_wire , x0x2x7_subscript1_share1_wire , x0x3x4_subscript1_share1_wire , x0x3x5_subscript1_share1_wire , x0x3x6_subscript1_share1_wire , x0x3x7_subscript1_share1_wire , x0x4x5_subscript1_share1_wire , x0x4x6_subscript1_share1_wire , x0x4x7_subscript1_share1_wire , x0x5x6_subscript1_share1_wire , x0x5x7_subscript1_share1_wire , x0x6x7_subscript1_share1_wire , x1x2x3_subscript1_share1_wire , x1x2x4_subscript1_share1_wire , x1x2x5_subscript1_share1_wire , x1x2x6_subscript1_share1_wire , x1x2x7_subscript1_share1_wire , x1x3x4_subscript1_share1_wire , x1x3x5_subscript1_share1_wire , x1x3x6_subscript1_share1_wire , x1x3x7_subscript1_share1_wire , x1x4x5_subscript1_share1_wire , x1x4x6_subscript1_share1_wire , x1x4x7_subscript1_share1_wire , x1x5x6_subscript1_share1_wire , x1x5x7_subscript1_share1_wire , x1x6x7_subscript1_share1_wire , x2x3x4_subscript1_share1_wire , x2x3x5_subscript1_share1_wire , x2x3x6_subscript1_share1_wire , x2x3x7_subscript1_share1_wire , x2x4x5_subscript1_share1_wire , x2x4x6_subscript1_share1_wire , x2x4x7_subscript1_share1_wire , x2x5x6_subscript1_share1_wire , x2x5x7_subscript1_share1_wire , x2x6x7_subscript1_share1_wire , x3x4x5_subscript1_share1_wire , x3x4x6_subscript1_share1_wire , x3x4x7_subscript1_share1_wire , x3x5x6_subscript1_share1_wire , x3x5x7_subscript1_share1_wire , x3x6x7_subscript1_share1_wire , x4x5x6_subscript1_share1_wire , x4x5x7_subscript1_share1_wire , x4x6x7_subscript1_share1_wire , x5x6x7_subscript1_share1_wire , x0x1x2x3_subscript1_share1_wire , x0x1x2x4_subscript1_share1_wire , x0x1x2x5_subscript1_share1_wire , x0x1x2x6_subscript1_share1_wire , x0x1x2x7_subscript1_share1_wire , x0x1x3x4_subscript1_share1_wire , x0x1x3x5_subscript1_share1_wire , x0x1x3x6_subscript1_share1_wire , x0x1x3x7_subscript1_share1_wire , x0x1x4x5_subscript1_share1_wire , x0x1x4x6_subscript1_share1_wire , x0x1x4x7_subscript1_share1_wire , x0x1x5x6_subscript1_share1_wire , x0x1x5x7_subscript1_share1_wire , x0x1x6x7_subscript1_share1_wire , x0x2x3x4_subscript1_share1_wire , x0x2x3x5_subscript1_share1_wire , x0x2x3x6_subscript1_share1_wire , x0x2x3x7_subscript1_share1_wire , x0x2x4x5_subscript1_share1_wire , x0x2x4x6_subscript1_share1_wire , x0x2x4x7_subscript1_share1_wire , x0x2x5x6_subscript1_share1_wire , x0x2x5x7_subscript1_share1_wire , x0x2x6x7_subscript1_share1_wire , x0x3x4x5_subscript1_share1_wire , x0x3x4x6_subscript1_share1_wire , x0x3x4x7_subscript1_share1_wire , x0x3x5x6_subscript1_share1_wire , x0x3x5x7_subscript1_share1_wire , x0x3x6x7_subscript1_share1_wire , x0x4x5x6_subscript1_share1_wire , x0x4x5x7_subscript1_share1_wire , x0x4x6x7_subscript1_share1_wire , x0x5x6x7_subscript1_share1_wire , x1x2x3x4_subscript1_share1_wire , x1x2x3x5_subscript1_share1_wire , x1x2x3x6_subscript1_share1_wire , x1x2x3x7_subscript1_share1_wire , x1x2x4x5_subscript1_share1_wire , x1x2x4x6_subscript1_share1_wire , x1x2x4x7_subscript1_share1_wire , x1x2x5x6_subscript1_share1_wire , x1x2x5x7_subscript1_share1_wire , x1x2x6x7_subscript1_share1_wire , x1x3x4x5_subscript1_share1_wire , x1x3x4x6_subscript1_share1_wire , x1x3x4x7_subscript1_share1_wire , x1x3x5x6_subscript1_share1_wire , x1x3x5x7_subscript1_share1_wire , x1x3x6x7_subscript1_share1_wire , x1x4x5x6_subscript1_share1_wire , x1x4x5x7_subscript1_share1_wire , x1x4x6x7_subscript1_share1_wire , x1x5x6x7_subscript1_share1_wire , x2x3x4x5_subscript1_share1_wire , x2x3x4x6_subscript1_share1_wire , x2x3x4x7_subscript1_share1_wire , x2x3x5x6_subscript1_share1_wire , x2x3x5x7_subscript1_share1_wire , x2x3x6x7_subscript1_share1_wire , x2x4x5x6_subscript1_share1_wire , x2x4x5x7_subscript1_share1_wire , x2x4x6x7_subscript1_share1_wire , x2x5x6x7_subscript1_share1_wire , x3x4x5x6_subscript1_share1_wire , x3x4x5x7_subscript1_share1_wire , x3x4x6x7_subscript1_share1_wire , x3x5x6x7_subscript1_share1_wire , x4x5x6x7_subscript1_share1_wire , x0x1x2x3x4_subscript1_share1_wire , x0x1x2x3x5_subscript1_share1_wire , x0x1x2x3x6_subscript1_share1_wire , x0x1x2x3x7_subscript1_share1_wire , x0x1x2x4x5_subscript1_share1_wire , x0x1x2x4x6_subscript1_share1_wire , x0x1x2x4x7_subscript1_share1_wire , x0x1x2x5x6_subscript1_share1_wire , x0x1x2x5x7_subscript1_share1_wire , x0x1x2x6x7_subscript1_share1_wire , x0x1x3x4x5_subscript1_share1_wire , x0x1x3x4x6_subscript1_share1_wire , x0x1x3x4x7_subscript1_share1_wire , x0x1x3x5x6_subscript1_share1_wire , x0x1x3x5x7_subscript1_share1_wire , x0x1x3x6x7_subscript1_share1_wire , x0x1x4x5x6_subscript1_share1_wire , x0x1x4x5x7_subscript1_share1_wire , x0x1x4x6x7_subscript1_share1_wire , x0x1x5x6x7_subscript1_share1_wire , x0x2x3x4x5_subscript1_share1_wire , x0x2x3x4x6_subscript1_share1_wire , x0x2x3x4x7_subscript1_share1_wire , x0x2x3x5x6_subscript1_share1_wire , x0x2x3x5x7_subscript1_share1_wire , x0x2x3x6x7_subscript1_share1_wire , x0x2x4x5x6_subscript1_share1_wire , x0x2x4x5x7_subscript1_share1_wire , x0x2x4x6x7_subscript1_share1_wire , x0x2x5x6x7_subscript1_share1_wire , x0x3x4x5x6_subscript1_share1_wire , x0x3x4x5x7_subscript1_share1_wire , x0x3x4x6x7_subscript1_share1_wire , x0x3x5x6x7_subscript1_share1_wire , x0x4x5x6x7_subscript1_share1_wire , x1x2x3x4x5_subscript1_share1_wire , x1x2x3x4x6_subscript1_share1_wire , x1x2x3x4x7_subscript1_share1_wire , x1x2x3x5x6_subscript1_share1_wire , x1x2x3x5x7_subscript1_share1_wire , x1x2x3x6x7_subscript1_share1_wire , x1x2x4x5x6_subscript1_share1_wire , x1x2x4x5x7_subscript1_share1_wire , x1x2x4x6x7_subscript1_share1_wire , x1x2x5x6x7_subscript1_share1_wire , x1x3x4x5x6_subscript1_share1_wire , x1x3x4x5x7_subscript1_share1_wire , x1x3x4x6x7_subscript1_share1_wire , x1x3x5x6x7_subscript1_share1_wire , x1x4x5x6x7_subscript1_share1_wire , x2x3x4x5x6_subscript1_share1_wire , x2x3x4x5x7_subscript1_share1_wire , x2x3x4x6x7_subscript1_share1_wire , x2x3x5x6x7_subscript1_share1_wire , x2x4x5x6x7_subscript1_share1_wire , x3x4x5x6x7_subscript1_share1_wire , x0x1x2x3x4x5_subscript1_share1_wire , x0x1x2x3x4x6_subscript1_share1_wire , x0x1x2x3x4x7_subscript1_share1_wire , x0x1x2x3x5x6_subscript1_share1_wire , x0x1x2x3x5x7_subscript1_share1_wire , x0x1x2x3x6x7_subscript1_share1_wire , x0x1x2x4x5x6_subscript1_share1_wire , x0x1x2x4x5x7_subscript1_share1_wire , x0x1x2x4x6x7_subscript1_share1_wire , x0x1x2x5x6x7_subscript1_share1_wire , x0x1x3x4x5x6_subscript1_share1_wire , x0x1x3x4x5x7_subscript1_share1_wire , x0x1x3x4x6x7_subscript1_share1_wire , x0x1x3x5x6x7_subscript1_share1_wire , x0x1x4x5x6x7_subscript1_share1_wire , x0x2x3x4x5x6_subscript1_share1_wire , x0x2x3x4x5x7_subscript1_share1_wire , x0x2x3x4x6x7_subscript1_share1_wire , x0x2x3x5x6x7_subscript1_share1_wire , x0x2x4x5x6x7_subscript1_share1_wire , x0x3x4x5x6x7_subscript1_share1_wire , x1x2x3x4x5x6_subscript1_share1_wire , x1x2x3x4x5x7_subscript1_share1_wire , x1x2x3x4x6x7_subscript1_share1_wire , x1x2x3x5x6x7_subscript1_share1_wire , x1x2x4x5x6x7_subscript1_share1_wire , x1x3x4x5x6x7_subscript1_share1_wire , x2x3x4x5x6x7_subscript1_share1_wire , x0x1x2x3x4x5x6_subscript1_share1_wire , x0x1x2x3x4x5x7_subscript1_share1_wire , x0x1x2x3x4x6x7_subscript1_share1_wire , x0x1x2x3x5x6x7_subscript1_share1_wire , x0x1x2x4x5x6x7_subscript1_share1_wire , x0x1x3x4x5x6x7_subscript1_share1_wire , x0x2x3x4x5x6x7_subscript1_share1_wire , x1x2x3x4x5x6x7_subscript1_share1_wire 
);

xor_AES_twofiftyfour xor_second_cycle_second_share(
    x0_subscript1_share2, x1_subscript1_share2, x2_subscript1_share2, x3_subscript1_share2, x4_subscript1_share2, x5_subscript1_share2, x6_subscript1_share2, x7_subscript1_share2 , x0x1_subscript1_share2 , x0x2_subscript1_share2 , x0x3_subscript1_share2 , x0x4_subscript1_share2 , x0x5_subscript1_share2 , x0x6_subscript1_share2 , x0x7_subscript1_share2 , x1x2_subscript1_share2 , x1x3_subscript1_share2 , x1x4_subscript1_share2 , x1x5_subscript1_share2 , x1x6_subscript1_share2 , x1x7_subscript1_share2 , x2x3_subscript1_share2 , x2x4_subscript1_share2 , x2x5_subscript1_share2 , x2x6_subscript1_share2 , x2x7_subscript1_share2 , x3x4_subscript1_share2 , x3x5_subscript1_share2 , x3x6_subscript1_share2 , x3x7_subscript1_share2 , x4x5_subscript1_share2 , x4x6_subscript1_share2 , x4x7_subscript1_share2 , x5x6_subscript1_share2 , x5x7_subscript1_share2 , x6x7_subscript1_share2 , x0x1x2_subscript1_share2 , x0x1x3_subscript1_share2 , x0x1x4_subscript1_share2 , x0x1x5_subscript1_share2 , x0x1x6_subscript1_share2 , x0x1x7_subscript1_share2 , x0x2x3_subscript1_share2 , x0x2x4_subscript1_share2 , x0x2x5_subscript1_share2 , x0x2x6_subscript1_share2 , x0x2x7_subscript1_share2 , x0x3x4_subscript1_share2 , x0x3x5_subscript1_share2 , x0x3x6_subscript1_share2 , x0x3x7_subscript1_share2 , x0x4x5_subscript1_share2 , x0x4x6_subscript1_share2 , x0x4x7_subscript1_share2 , x0x5x6_subscript1_share2 , x0x5x7_subscript1_share2 , x0x6x7_subscript1_share2 , x1x2x3_subscript1_share2 , x1x2x4_subscript1_share2 , x1x2x5_subscript1_share2 , x1x2x6_subscript1_share2 , x1x2x7_subscript1_share2 , x1x3x4_subscript1_share2 , x1x3x5_subscript1_share2 , x1x3x6_subscript1_share2 , x1x3x7_subscript1_share2 , x1x4x5_subscript1_share2 , x1x4x6_subscript1_share2 , x1x4x7_subscript1_share2 , x1x5x6_subscript1_share2 , x1x5x7_subscript1_share2 , x1x6x7_subscript1_share2 , x2x3x4_subscript1_share2 , x2x3x5_subscript1_share2 , x2x3x6_subscript1_share2 , x2x3x7_subscript1_share2 , x2x4x5_subscript1_share2 , x2x4x6_subscript1_share2 , x2x4x7_subscript1_share2 , x2x5x6_subscript1_share2 , x2x5x7_subscript1_share2 , x2x6x7_subscript1_share2 , x3x4x5_subscript1_share2 , x3x4x6_subscript1_share2 , x3x4x7_subscript1_share2 , x3x5x6_subscript1_share2 , x3x5x7_subscript1_share2 , x3x6x7_subscript1_share2 , x4x5x6_subscript1_share2 , x4x5x7_subscript1_share2 , x4x6x7_subscript1_share2 , x5x6x7_subscript1_share2 , x0x1x2x3_subscript1_share2 , x0x1x2x4_subscript1_share2 , x0x1x2x5_subscript1_share2 , x0x1x2x6_subscript1_share2 , x0x1x2x7_subscript1_share2 , x0x1x3x4_subscript1_share2 , x0x1x3x5_subscript1_share2 , x0x1x3x6_subscript1_share2 , x0x1x3x7_subscript1_share2 , x0x1x4x5_subscript1_share2 , x0x1x4x6_subscript1_share2 , x0x1x4x7_subscript1_share2 , x0x1x5x6_subscript1_share2 , x0x1x5x7_subscript1_share2 , x0x1x6x7_subscript1_share2 , x0x2x3x4_subscript1_share2 , x0x2x3x5_subscript1_share2 , x0x2x3x6_subscript1_share2 , x0x2x3x7_subscript1_share2 , x0x2x4x5_subscript1_share2 , x0x2x4x6_subscript1_share2 , x0x2x4x7_subscript1_share2 , x0x2x5x6_subscript1_share2 , x0x2x5x7_subscript1_share2 , x0x2x6x7_subscript1_share2 , x0x3x4x5_subscript1_share2 , x0x3x4x6_subscript1_share2 , x0x3x4x7_subscript1_share2 , x0x3x5x6_subscript1_share2 , x0x3x5x7_subscript1_share2 , x0x3x6x7_subscript1_share2 , x0x4x5x6_subscript1_share2 , x0x4x5x7_subscript1_share2 , x0x4x6x7_subscript1_share2 , x0x5x6x7_subscript1_share2 , x1x2x3x4_subscript1_share2 , x1x2x3x5_subscript1_share2 , x1x2x3x6_subscript1_share2 , x1x2x3x7_subscript1_share2 , x1x2x4x5_subscript1_share2 , x1x2x4x6_subscript1_share2 , x1x2x4x7_subscript1_share2 , x1x2x5x6_subscript1_share2 , x1x2x5x7_subscript1_share2 , x1x2x6x7_subscript1_share2 , x1x3x4x5_subscript1_share2 , x1x3x4x6_subscript1_share2 , x1x3x4x7_subscript1_share2 , x1x3x5x6_subscript1_share2 , x1x3x5x7_subscript1_share2 , x1x3x6x7_subscript1_share2 , x1x4x5x6_subscript1_share2 , x1x4x5x7_subscript1_share2 , x1x4x6x7_subscript1_share2 , x1x5x6x7_subscript1_share2 , x2x3x4x5_subscript1_share2 , x2x3x4x6_subscript1_share2 , x2x3x4x7_subscript1_share2 , x2x3x5x6_subscript1_share2 , x2x3x5x7_subscript1_share2 , x2x3x6x7_subscript1_share2 , x2x4x5x6_subscript1_share2 , x2x4x5x7_subscript1_share2 , x2x4x6x7_subscript1_share2 , x2x5x6x7_subscript1_share2 , x3x4x5x6_subscript1_share2 , x3x4x5x7_subscript1_share2 , x3x4x6x7_subscript1_share2 , x3x5x6x7_subscript1_share2 , x4x5x6x7_subscript1_share2 , x0x1x2x3x4_subscript1_share2 , x0x1x2x3x5_subscript1_share2 , x0x1x2x3x6_subscript1_share2 , x0x1x2x3x7_subscript1_share2 , x0x1x2x4x5_subscript1_share2 , x0x1x2x4x6_subscript1_share2 , x0x1x2x4x7_subscript1_share2 , x0x1x2x5x6_subscript1_share2 , x0x1x2x5x7_subscript1_share2 , x0x1x2x6x7_subscript1_share2 , x0x1x3x4x5_subscript1_share2 , x0x1x3x4x6_subscript1_share2 , x0x1x3x4x7_subscript1_share2 , x0x1x3x5x6_subscript1_share2 , x0x1x3x5x7_subscript1_share2 , x0x1x3x6x7_subscript1_share2 , x0x1x4x5x6_subscript1_share2 , x0x1x4x5x7_subscript1_share2 , x0x1x4x6x7_subscript1_share2 , x0x1x5x6x7_subscript1_share2 , x0x2x3x4x5_subscript1_share2 , x0x2x3x4x6_subscript1_share2 , x0x2x3x4x7_subscript1_share2 , x0x2x3x5x6_subscript1_share2 , x0x2x3x5x7_subscript1_share2 , x0x2x3x6x7_subscript1_share2 , x0x2x4x5x6_subscript1_share2 , x0x2x4x5x7_subscript1_share2 , x0x2x4x6x7_subscript1_share2 , x0x2x5x6x7_subscript1_share2 , x0x3x4x5x6_subscript1_share2 , x0x3x4x5x7_subscript1_share2 , x0x3x4x6x7_subscript1_share2 , x0x3x5x6x7_subscript1_share2 , x0x4x5x6x7_subscript1_share2 , x1x2x3x4x5_subscript1_share2 , x1x2x3x4x6_subscript1_share2 , x1x2x3x4x7_subscript1_share2 , x1x2x3x5x6_subscript1_share2 , x1x2x3x5x7_subscript1_share2 , x1x2x3x6x7_subscript1_share2 , x1x2x4x5x6_subscript1_share2 , x1x2x4x5x7_subscript1_share2 , x1x2x4x6x7_subscript1_share2 , x1x2x5x6x7_subscript1_share2 , x1x3x4x5x6_subscript1_share2 , x1x3x4x5x7_subscript1_share2 , x1x3x4x6x7_subscript1_share2 , x1x3x5x6x7_subscript1_share2 , x1x4x5x6x7_subscript1_share2 , x2x3x4x5x6_subscript1_share2 , x2x3x4x5x7_subscript1_share2 , x2x3x4x6x7_subscript1_share2 , x2x3x5x6x7_subscript1_share2 , x2x4x5x6x7_subscript1_share2 , x3x4x5x6x7_subscript1_share2 , x0x1x2x3x4x5_subscript1_share2 , x0x1x2x3x4x6_subscript1_share2 , x0x1x2x3x4x7_subscript1_share2 , x0x1x2x3x5x6_subscript1_share2 , x0x1x2x3x5x7_subscript1_share2 , x0x1x2x3x6x7_subscript1_share2 , x0x1x2x4x5x6_subscript1_share2 , x0x1x2x4x5x7_subscript1_share2 , x0x1x2x4x6x7_subscript1_share2 , x0x1x2x5x6x7_subscript1_share2 , x0x1x3x4x5x6_subscript1_share2 , x0x1x3x4x5x7_subscript1_share2 , x0x1x3x4x6x7_subscript1_share2 , x0x1x3x5x6x7_subscript1_share2 , x0x1x4x5x6x7_subscript1_share2 , x0x2x3x4x5x6_subscript1_share2 , x0x2x3x4x5x7_subscript1_share2 , x0x2x3x4x6x7_subscript1_share2 , x0x2x3x5x6x7_subscript1_share2 , x0x2x4x5x6x7_subscript1_share2 , x0x3x4x5x6x7_subscript1_share2 , x1x2x3x4x5x6_subscript1_share2 , x1x2x3x4x5x7_subscript1_share2 , x1x2x3x4x6x7_subscript1_share2 , x1x2x3x5x6x7_subscript1_share2 , x1x2x4x5x6x7_subscript1_share2 , x1x3x4x5x6x7_subscript1_share2 , x2x3x4x5x6x7_subscript1_share2 , x0x1x2x3x4x5x6_subscript1_share2 , x0x1x2x3x4x5x7_subscript1_share2 , x0x1x2x3x4x6x7_subscript1_share2 , x0x1x2x3x5x6x7_subscript1_share2 , x0x1x2x4x5x6x7_subscript1_share2 , x0x1x3x4x5x6x7_subscript1_share2 , x0x2x3x4x5x6x7_subscript1_share2 , x1x2x3x4x5x6x7_subscript1_share2 ,
    rand_second_cycle_b[1] ,rand_second_cycle_b[2] ,rand_second_cycle_b[3] ,rand_second_cycle_b[4] ,rand_second_cycle_b[5] ,rand_second_cycle_b[6] ,rand_second_cycle_b[7] ,rand_second_cycle_b[8] ,rand_second_cycle_b[9] ,rand_second_cycle_b[10] ,rand_second_cycle_b[11] ,rand_second_cycle_b[12] ,rand_second_cycle_b[13] ,rand_second_cycle_b[14] ,rand_second_cycle_b[15] ,rand_second_cycle_b[16] ,rand_second_cycle_b[17] ,rand_second_cycle_b[18] ,rand_second_cycle_b[19] ,rand_second_cycle_b[20] ,rand_second_cycle_b[21] ,rand_second_cycle_b[22] ,rand_second_cycle_b[23] ,rand_second_cycle_b[24] ,rand_second_cycle_b[25] ,rand_second_cycle_b[26] ,rand_second_cycle_b[27] ,rand_second_cycle_b[28] ,rand_second_cycle_b[29] ,rand_second_cycle_b[30] ,rand_second_cycle_b[31] ,rand_second_cycle_b[32] ,rand_second_cycle_b[33] ,rand_second_cycle_b[34] ,rand_second_cycle_b[35] ,rand_second_cycle_b[36] ,rand_second_cycle_b[37] ,rand_second_cycle_b[38] ,rand_second_cycle_b[39] ,rand_second_cycle_b[40] ,rand_second_cycle_b[41] ,rand_second_cycle_b[42] ,rand_second_cycle_b[43] ,rand_second_cycle_b[44] ,rand_second_cycle_b[45] ,rand_second_cycle_b[46] ,rand_second_cycle_b[47] ,rand_second_cycle_b[48] ,rand_second_cycle_b[49] ,rand_second_cycle_b[50] ,rand_second_cycle_b[51] ,rand_second_cycle_b[52] ,rand_second_cycle_b[53] ,rand_second_cycle_b[54] ,rand_second_cycle_b[55] ,rand_second_cycle_b[56] ,rand_second_cycle_b[57] ,rand_second_cycle_b[58] ,rand_second_cycle_b[59] ,rand_second_cycle_b[60] ,rand_second_cycle_b[61] ,rand_second_cycle_b[62] ,rand_second_cycle_b[63] ,rand_second_cycle_b[64] ,rand_second_cycle_b[65] ,rand_second_cycle_b[66] ,rand_second_cycle_b[67] ,rand_second_cycle_b[68] ,rand_second_cycle_b[69] ,rand_second_cycle_b[70] ,rand_second_cycle_b[71] ,rand_second_cycle_b[72] ,rand_second_cycle_b[73] ,rand_second_cycle_b[74] ,rand_second_cycle_b[75] ,rand_second_cycle_b[76] ,rand_second_cycle_b[77] ,rand_second_cycle_b[78] ,rand_second_cycle_b[79] ,rand_second_cycle_b[80] ,rand_second_cycle_b[81] ,rand_second_cycle_b[82] ,rand_second_cycle_b[83] ,rand_second_cycle_b[84] ,rand_second_cycle_b[85] ,rand_second_cycle_b[86] ,rand_second_cycle_b[87] ,rand_second_cycle_b[88] ,rand_second_cycle_b[89] ,rand_second_cycle_b[90] ,rand_second_cycle_b[91] ,rand_second_cycle_b[92] ,rand_second_cycle_b[93] ,rand_second_cycle_b[94] ,rand_second_cycle_b[95] ,rand_second_cycle_b[96] ,rand_second_cycle_b[97] ,rand_second_cycle_b[98] ,rand_second_cycle_b[99] ,rand_second_cycle_b[100] ,rand_second_cycle_b[101] ,rand_second_cycle_b[102] ,rand_second_cycle_b[103] ,rand_second_cycle_b[104] ,rand_second_cycle_b[105] ,rand_second_cycle_b[106] ,rand_second_cycle_b[107] ,rand_second_cycle_b[108] ,rand_second_cycle_b[109] ,rand_second_cycle_b[110] ,rand_second_cycle_b[111] ,rand_second_cycle_b[112] ,rand_second_cycle_b[113] ,rand_second_cycle_b[114] ,rand_second_cycle_b[115] ,rand_second_cycle_b[116] ,rand_second_cycle_b[117] ,rand_second_cycle_b[118] ,rand_second_cycle_b[119] ,rand_second_cycle_b[120] ,rand_second_cycle_b[121] ,rand_second_cycle_b[122] ,rand_second_cycle_b[123] ,rand_second_cycle_b[124] ,rand_second_cycle_b[125] ,rand_second_cycle_b[126] ,rand_second_cycle_b[127] ,rand_second_cycle_b[128] ,rand_second_cycle_b[129] ,rand_second_cycle_b[130] ,rand_second_cycle_b[131] ,rand_second_cycle_b[132] ,rand_second_cycle_b[133] ,rand_second_cycle_b[134] ,rand_second_cycle_b[135] ,rand_second_cycle_b[136] ,rand_second_cycle_b[137] ,rand_second_cycle_b[138] ,rand_second_cycle_b[139] ,rand_second_cycle_b[140] ,rand_second_cycle_b[141] ,rand_second_cycle_b[142] ,rand_second_cycle_b[143] ,rand_second_cycle_b[144] ,rand_second_cycle_b[145] ,rand_second_cycle_b[146] ,rand_second_cycle_b[147] ,rand_second_cycle_b[148] ,rand_second_cycle_b[149] ,rand_second_cycle_b[150] ,rand_second_cycle_b[151] ,rand_second_cycle_b[152] ,rand_second_cycle_b[153] ,rand_second_cycle_b[154] ,rand_second_cycle_b[155] ,rand_second_cycle_b[156] ,rand_second_cycle_b[157] ,rand_second_cycle_b[158] ,rand_second_cycle_b[159] ,rand_second_cycle_b[160] ,rand_second_cycle_b[161] ,rand_second_cycle_b[162] ,rand_second_cycle_b[163] ,rand_second_cycle_b[164] ,rand_second_cycle_b[165] ,rand_second_cycle_b[166] ,rand_second_cycle_b[167] ,rand_second_cycle_b[168] ,rand_second_cycle_b[169] ,rand_second_cycle_b[170] ,rand_second_cycle_b[171] ,rand_second_cycle_b[172] ,rand_second_cycle_b[173] ,rand_second_cycle_b[174] ,rand_second_cycle_b[175] ,rand_second_cycle_b[176] ,rand_second_cycle_b[177] ,rand_second_cycle_b[178] ,rand_second_cycle_b[179] ,rand_second_cycle_b[180] ,rand_second_cycle_b[181] ,rand_second_cycle_b[182] ,rand_second_cycle_b[183] ,rand_second_cycle_b[184] ,rand_second_cycle_b[185] ,rand_second_cycle_b[186] ,rand_second_cycle_b[187] ,rand_second_cycle_b[188] ,rand_second_cycle_b[189] ,rand_second_cycle_b[190] ,rand_second_cycle_b[191] ,rand_second_cycle_b[192] ,rand_second_cycle_b[193] ,rand_second_cycle_b[194] ,rand_second_cycle_b[195] ,rand_second_cycle_b[196] ,rand_second_cycle_b[197] ,rand_second_cycle_b[198] ,rand_second_cycle_b[199] ,rand_second_cycle_b[200] ,rand_second_cycle_b[201] ,rand_second_cycle_b[202] ,rand_second_cycle_b[203] ,rand_second_cycle_b[204] ,rand_second_cycle_b[205] ,rand_second_cycle_b[206] ,rand_second_cycle_b[207] ,rand_second_cycle_b[208] ,rand_second_cycle_b[209] ,rand_second_cycle_b[210] ,rand_second_cycle_b[211] ,rand_second_cycle_b[212] ,rand_second_cycle_b[213] ,rand_second_cycle_b[214] ,rand_second_cycle_b[215] ,rand_second_cycle_b[216] ,rand_second_cycle_b[217] ,rand_second_cycle_b[218] ,rand_second_cycle_b[219] ,rand_second_cycle_b[220] ,rand_second_cycle_b[221] ,rand_second_cycle_b[222] ,rand_second_cycle_b[223] ,rand_second_cycle_b[224] ,rand_second_cycle_b[225] ,rand_second_cycle_b[226] ,rand_second_cycle_b[227] ,rand_second_cycle_b[228] ,rand_second_cycle_b[229] ,rand_second_cycle_b[230] ,rand_second_cycle_b[231] ,rand_second_cycle_b[232] ,rand_second_cycle_b[233] ,rand_second_cycle_b[234] ,rand_second_cycle_b[235] ,rand_second_cycle_b[236] ,rand_second_cycle_b[237] ,rand_second_cycle_b[238] ,rand_second_cycle_b[239] ,rand_second_cycle_b[240] ,rand_second_cycle_b[241] ,rand_second_cycle_b[242] ,rand_second_cycle_b[243] ,rand_second_cycle_b[244] ,rand_second_cycle_b[245] ,rand_second_cycle_b[246] ,rand_second_cycle_b[247] ,rand_second_cycle_b[248] ,rand_second_cycle_b[249] ,rand_second_cycle_b[250] ,rand_second_cycle_b[251] ,rand_second_cycle_b[252] ,rand_second_cycle_b[253] ,rand_second_cycle_b[254] ,
    x0_subscript1_share2_wire, x1_subscript1_share2_wire, x2_subscript1_share2_wire, x3_subscript1_share2_wire, x4_subscript1_share2_wire, x5_subscript1_share2_wire, x6_subscript1_share2_wire, x7_subscript1_share2_wire , x0x1_subscript1_share2_wire , x0x2_subscript1_share2_wire , x0x3_subscript1_share2_wire , x0x4_subscript1_share2_wire , x0x5_subscript1_share2_wire , x0x6_subscript1_share2_wire , x0x7_subscript1_share2_wire , x1x2_subscript1_share2_wire , x1x3_subscript1_share2_wire , x1x4_subscript1_share2_wire , x1x5_subscript1_share2_wire , x1x6_subscript1_share2_wire , x1x7_subscript1_share2_wire , x2x3_subscript1_share2_wire , x2x4_subscript1_share2_wire , x2x5_subscript1_share2_wire , x2x6_subscript1_share2_wire , x2x7_subscript1_share2_wire , x3x4_subscript1_share2_wire , x3x5_subscript1_share2_wire , x3x6_subscript1_share2_wire , x3x7_subscript1_share2_wire , x4x5_subscript1_share2_wire , x4x6_subscript1_share2_wire , x4x7_subscript1_share2_wire , x5x6_subscript1_share2_wire , x5x7_subscript1_share2_wire , x6x7_subscript1_share2_wire , x0x1x2_subscript1_share2_wire , x0x1x3_subscript1_share2_wire , x0x1x4_subscript1_share2_wire , x0x1x5_subscript1_share2_wire , x0x1x6_subscript1_share2_wire , x0x1x7_subscript1_share2_wire , x0x2x3_subscript1_share2_wire , x0x2x4_subscript1_share2_wire , x0x2x5_subscript1_share2_wire , x0x2x6_subscript1_share2_wire , x0x2x7_subscript1_share2_wire , x0x3x4_subscript1_share2_wire , x0x3x5_subscript1_share2_wire , x0x3x6_subscript1_share2_wire , x0x3x7_subscript1_share2_wire , x0x4x5_subscript1_share2_wire , x0x4x6_subscript1_share2_wire , x0x4x7_subscript1_share2_wire , x0x5x6_subscript1_share2_wire , x0x5x7_subscript1_share2_wire , x0x6x7_subscript1_share2_wire , x1x2x3_subscript1_share2_wire , x1x2x4_subscript1_share2_wire , x1x2x5_subscript1_share2_wire , x1x2x6_subscript1_share2_wire , x1x2x7_subscript1_share2_wire , x1x3x4_subscript1_share2_wire , x1x3x5_subscript1_share2_wire , x1x3x6_subscript1_share2_wire , x1x3x7_subscript1_share2_wire , x1x4x5_subscript1_share2_wire , x1x4x6_subscript1_share2_wire , x1x4x7_subscript1_share2_wire , x1x5x6_subscript1_share2_wire , x1x5x7_subscript1_share2_wire , x1x6x7_subscript1_share2_wire , x2x3x4_subscript1_share2_wire , x2x3x5_subscript1_share2_wire , x2x3x6_subscript1_share2_wire , x2x3x7_subscript1_share2_wire , x2x4x5_subscript1_share2_wire , x2x4x6_subscript1_share2_wire , x2x4x7_subscript1_share2_wire , x2x5x6_subscript1_share2_wire , x2x5x7_subscript1_share2_wire , x2x6x7_subscript1_share2_wire , x3x4x5_subscript1_share2_wire , x3x4x6_subscript1_share2_wire , x3x4x7_subscript1_share2_wire , x3x5x6_subscript1_share2_wire , x3x5x7_subscript1_share2_wire , x3x6x7_subscript1_share2_wire , x4x5x6_subscript1_share2_wire , x4x5x7_subscript1_share2_wire , x4x6x7_subscript1_share2_wire , x5x6x7_subscript1_share2_wire , x0x1x2x3_subscript1_share2_wire , x0x1x2x4_subscript1_share2_wire , x0x1x2x5_subscript1_share2_wire , x0x1x2x6_subscript1_share2_wire , x0x1x2x7_subscript1_share2_wire , x0x1x3x4_subscript1_share2_wire , x0x1x3x5_subscript1_share2_wire , x0x1x3x6_subscript1_share2_wire , x0x1x3x7_subscript1_share2_wire , x0x1x4x5_subscript1_share2_wire , x0x1x4x6_subscript1_share2_wire , x0x1x4x7_subscript1_share2_wire , x0x1x5x6_subscript1_share2_wire , x0x1x5x7_subscript1_share2_wire , x0x1x6x7_subscript1_share2_wire , x0x2x3x4_subscript1_share2_wire , x0x2x3x5_subscript1_share2_wire , x0x2x3x6_subscript1_share2_wire , x0x2x3x7_subscript1_share2_wire , x0x2x4x5_subscript1_share2_wire , x0x2x4x6_subscript1_share2_wire , x0x2x4x7_subscript1_share2_wire , x0x2x5x6_subscript1_share2_wire , x0x2x5x7_subscript1_share2_wire , x0x2x6x7_subscript1_share2_wire , x0x3x4x5_subscript1_share2_wire , x0x3x4x6_subscript1_share2_wire , x0x3x4x7_subscript1_share2_wire , x0x3x5x6_subscript1_share2_wire , x0x3x5x7_subscript1_share2_wire , x0x3x6x7_subscript1_share2_wire , x0x4x5x6_subscript1_share2_wire , x0x4x5x7_subscript1_share2_wire , x0x4x6x7_subscript1_share2_wire , x0x5x6x7_subscript1_share2_wire , x1x2x3x4_subscript1_share2_wire , x1x2x3x5_subscript1_share2_wire , x1x2x3x6_subscript1_share2_wire , x1x2x3x7_subscript1_share2_wire , x1x2x4x5_subscript1_share2_wire , x1x2x4x6_subscript1_share2_wire , x1x2x4x7_subscript1_share2_wire , x1x2x5x6_subscript1_share2_wire , x1x2x5x7_subscript1_share2_wire , x1x2x6x7_subscript1_share2_wire , x1x3x4x5_subscript1_share2_wire , x1x3x4x6_subscript1_share2_wire , x1x3x4x7_subscript1_share2_wire , x1x3x5x6_subscript1_share2_wire , x1x3x5x7_subscript1_share2_wire , x1x3x6x7_subscript1_share2_wire , x1x4x5x6_subscript1_share2_wire , x1x4x5x7_subscript1_share2_wire , x1x4x6x7_subscript1_share2_wire , x1x5x6x7_subscript1_share2_wire , x2x3x4x5_subscript1_share2_wire , x2x3x4x6_subscript1_share2_wire , x2x3x4x7_subscript1_share2_wire , x2x3x5x6_subscript1_share2_wire , x2x3x5x7_subscript1_share2_wire , x2x3x6x7_subscript1_share2_wire , x2x4x5x6_subscript1_share2_wire , x2x4x5x7_subscript1_share2_wire , x2x4x6x7_subscript1_share2_wire , x2x5x6x7_subscript1_share2_wire , x3x4x5x6_subscript1_share2_wire , x3x4x5x7_subscript1_share2_wire , x3x4x6x7_subscript1_share2_wire , x3x5x6x7_subscript1_share2_wire , x4x5x6x7_subscript1_share2_wire , x0x1x2x3x4_subscript1_share2_wire , x0x1x2x3x5_subscript1_share2_wire , x0x1x2x3x6_subscript1_share2_wire , x0x1x2x3x7_subscript1_share2_wire , x0x1x2x4x5_subscript1_share2_wire , x0x1x2x4x6_subscript1_share2_wire , x0x1x2x4x7_subscript1_share2_wire , x0x1x2x5x6_subscript1_share2_wire , x0x1x2x5x7_subscript1_share2_wire , x0x1x2x6x7_subscript1_share2_wire , x0x1x3x4x5_subscript1_share2_wire , x0x1x3x4x6_subscript1_share2_wire , x0x1x3x4x7_subscript1_share2_wire , x0x1x3x5x6_subscript1_share2_wire , x0x1x3x5x7_subscript1_share2_wire , x0x1x3x6x7_subscript1_share2_wire , x0x1x4x5x6_subscript1_share2_wire , x0x1x4x5x7_subscript1_share2_wire , x0x1x4x6x7_subscript1_share2_wire , x0x1x5x6x7_subscript1_share2_wire , x0x2x3x4x5_subscript1_share2_wire , x0x2x3x4x6_subscript1_share2_wire , x0x2x3x4x7_subscript1_share2_wire , x0x2x3x5x6_subscript1_share2_wire , x0x2x3x5x7_subscript1_share2_wire , x0x2x3x6x7_subscript1_share2_wire , x0x2x4x5x6_subscript1_share2_wire , x0x2x4x5x7_subscript1_share2_wire , x0x2x4x6x7_subscript1_share2_wire , x0x2x5x6x7_subscript1_share2_wire , x0x3x4x5x6_subscript1_share2_wire , x0x3x4x5x7_subscript1_share2_wire , x0x3x4x6x7_subscript1_share2_wire , x0x3x5x6x7_subscript1_share2_wire , x0x4x5x6x7_subscript1_share2_wire , x1x2x3x4x5_subscript1_share2_wire , x1x2x3x4x6_subscript1_share2_wire , x1x2x3x4x7_subscript1_share2_wire , x1x2x3x5x6_subscript1_share2_wire , x1x2x3x5x7_subscript1_share2_wire , x1x2x3x6x7_subscript1_share2_wire , x1x2x4x5x6_subscript1_share2_wire , x1x2x4x5x7_subscript1_share2_wire , x1x2x4x6x7_subscript1_share2_wire , x1x2x5x6x7_subscript1_share2_wire , x1x3x4x5x6_subscript1_share2_wire , x1x3x4x5x7_subscript1_share2_wire , x1x3x4x6x7_subscript1_share2_wire , x1x3x5x6x7_subscript1_share2_wire , x1x4x5x6x7_subscript1_share2_wire , x2x3x4x5x6_subscript1_share2_wire , x2x3x4x5x7_subscript1_share2_wire , x2x3x4x6x7_subscript1_share2_wire , x2x3x5x6x7_subscript1_share2_wire , x2x4x5x6x7_subscript1_share2_wire , x3x4x5x6x7_subscript1_share2_wire , x0x1x2x3x4x5_subscript1_share2_wire , x0x1x2x3x4x6_subscript1_share2_wire , x0x1x2x3x4x7_subscript1_share2_wire , x0x1x2x3x5x6_subscript1_share2_wire , x0x1x2x3x5x7_subscript1_share2_wire , x0x1x2x3x6x7_subscript1_share2_wire , x0x1x2x4x5x6_subscript1_share2_wire , x0x1x2x4x5x7_subscript1_share2_wire , x0x1x2x4x6x7_subscript1_share2_wire , x0x1x2x5x6x7_subscript1_share2_wire , x0x1x3x4x5x6_subscript1_share2_wire , x0x1x3x4x5x7_subscript1_share2_wire , x0x1x3x4x6x7_subscript1_share2_wire , x0x1x3x5x6x7_subscript1_share2_wire , x0x1x4x5x6x7_subscript1_share2_wire , x0x2x3x4x5x6_subscript1_share2_wire , x0x2x3x4x5x7_subscript1_share2_wire , x0x2x3x4x6x7_subscript1_share2_wire , x0x2x3x5x6x7_subscript1_share2_wire , x0x2x4x5x6x7_subscript1_share2_wire , x0x3x4x5x6x7_subscript1_share2_wire , x1x2x3x4x5x6_subscript1_share2_wire , x1x2x3x4x5x7_subscript1_share2_wire , x1x2x3x4x6x7_subscript1_share2_wire , x1x2x3x5x6x7_subscript1_share2_wire , x1x2x4x5x6x7_subscript1_share2_wire , x1x3x4x5x6x7_subscript1_share2_wire , x2x3x4x5x6x7_subscript1_share2_wire , x0x1x2x3x4x5x6_subscript1_share2_wire , x0x1x2x3x4x5x7_subscript1_share2_wire , x0x1x2x3x4x6x7_subscript1_share2_wire , x0x1x2x3x5x6x7_subscript1_share2_wire , x0x1x2x4x5x6x7_subscript1_share2_wire , x0x1x3x4x5x6x7_subscript1_share2_wire , x0x2x3x4x5x6x7_subscript1_share2_wire , x1x2x3x4x5x6x7_subscript1_share2_wire 
);

xor_AES_twofiftyfour xor_second_cycle_third_share(
    rand_second_cycle_a[1] ,rand_second_cycle_a[2] ,rand_second_cycle_a[3] ,rand_second_cycle_a[4] ,rand_second_cycle_a[5] ,rand_second_cycle_a[6] ,rand_second_cycle_a[7] ,rand_second_cycle_a[8] ,rand_second_cycle_a[9] ,rand_second_cycle_a[10] ,rand_second_cycle_a[11] ,rand_second_cycle_a[12] ,rand_second_cycle_a[13] ,rand_second_cycle_a[14] ,rand_second_cycle_a[15] ,rand_second_cycle_a[16] ,rand_second_cycle_a[17] ,rand_second_cycle_a[18] ,rand_second_cycle_a[19] ,rand_second_cycle_a[20] ,rand_second_cycle_a[21] ,rand_second_cycle_a[22] ,rand_second_cycle_a[23] ,rand_second_cycle_a[24] ,rand_second_cycle_a[25] ,rand_second_cycle_a[26] ,rand_second_cycle_a[27] ,rand_second_cycle_a[28] ,rand_second_cycle_a[29] ,rand_second_cycle_a[30] ,rand_second_cycle_a[31] ,rand_second_cycle_a[32] ,rand_second_cycle_a[33] ,rand_second_cycle_a[34] ,rand_second_cycle_a[35] ,rand_second_cycle_a[36] ,rand_second_cycle_a[37] ,rand_second_cycle_a[38] ,rand_second_cycle_a[39] ,rand_second_cycle_a[40] ,rand_second_cycle_a[41] ,rand_second_cycle_a[42] ,rand_second_cycle_a[43] ,rand_second_cycle_a[44] ,rand_second_cycle_a[45] ,rand_second_cycle_a[46] ,rand_second_cycle_a[47] ,rand_second_cycle_a[48] ,rand_second_cycle_a[49] ,rand_second_cycle_a[50] ,rand_second_cycle_a[51] ,rand_second_cycle_a[52] ,rand_second_cycle_a[53] ,rand_second_cycle_a[54] ,rand_second_cycle_a[55] ,rand_second_cycle_a[56] ,rand_second_cycle_a[57] ,rand_second_cycle_a[58] ,rand_second_cycle_a[59] ,rand_second_cycle_a[60] ,rand_second_cycle_a[61] ,rand_second_cycle_a[62] ,rand_second_cycle_a[63] ,rand_second_cycle_a[64] ,rand_second_cycle_a[65] ,rand_second_cycle_a[66] ,rand_second_cycle_a[67] ,rand_second_cycle_a[68] ,rand_second_cycle_a[69] ,rand_second_cycle_a[70] ,rand_second_cycle_a[71] ,rand_second_cycle_a[72] ,rand_second_cycle_a[73] ,rand_second_cycle_a[74] ,rand_second_cycle_a[75] ,rand_second_cycle_a[76] ,rand_second_cycle_a[77] ,rand_second_cycle_a[78] ,rand_second_cycle_a[79] ,rand_second_cycle_a[80] ,rand_second_cycle_a[81] ,rand_second_cycle_a[82] ,rand_second_cycle_a[83] ,rand_second_cycle_a[84] ,rand_second_cycle_a[85] ,rand_second_cycle_a[86] ,rand_second_cycle_a[87] ,rand_second_cycle_a[88] ,rand_second_cycle_a[89] ,rand_second_cycle_a[90] ,rand_second_cycle_a[91] ,rand_second_cycle_a[92] ,rand_second_cycle_a[93] ,rand_second_cycle_a[94] ,rand_second_cycle_a[95] ,rand_second_cycle_a[96] ,rand_second_cycle_a[97] ,rand_second_cycle_a[98] ,rand_second_cycle_a[99] ,rand_second_cycle_a[100] ,rand_second_cycle_a[101] ,rand_second_cycle_a[102] ,rand_second_cycle_a[103] ,rand_second_cycle_a[104] ,rand_second_cycle_a[105] ,rand_second_cycle_a[106] ,rand_second_cycle_a[107] ,rand_second_cycle_a[108] ,rand_second_cycle_a[109] ,rand_second_cycle_a[110] ,rand_second_cycle_a[111] ,rand_second_cycle_a[112] ,rand_second_cycle_a[113] ,rand_second_cycle_a[114] ,rand_second_cycle_a[115] ,rand_second_cycle_a[116] ,rand_second_cycle_a[117] ,rand_second_cycle_a[118] ,rand_second_cycle_a[119] ,rand_second_cycle_a[120] ,rand_second_cycle_a[121] ,rand_second_cycle_a[122] ,rand_second_cycle_a[123] ,rand_second_cycle_a[124] ,rand_second_cycle_a[125] ,rand_second_cycle_a[126] ,rand_second_cycle_a[127] ,rand_second_cycle_a[128] ,rand_second_cycle_a[129] ,rand_second_cycle_a[130] ,rand_second_cycle_a[131] ,rand_second_cycle_a[132] ,rand_second_cycle_a[133] ,rand_second_cycle_a[134] ,rand_second_cycle_a[135] ,rand_second_cycle_a[136] ,rand_second_cycle_a[137] ,rand_second_cycle_a[138] ,rand_second_cycle_a[139] ,rand_second_cycle_a[140] ,rand_second_cycle_a[141] ,rand_second_cycle_a[142] ,rand_second_cycle_a[143] ,rand_second_cycle_a[144] ,rand_second_cycle_a[145] ,rand_second_cycle_a[146] ,rand_second_cycle_a[147] ,rand_second_cycle_a[148] ,rand_second_cycle_a[149] ,rand_second_cycle_a[150] ,rand_second_cycle_a[151] ,rand_second_cycle_a[152] ,rand_second_cycle_a[153] ,rand_second_cycle_a[154] ,rand_second_cycle_a[155] ,rand_second_cycle_a[156] ,rand_second_cycle_a[157] ,rand_second_cycle_a[158] ,rand_second_cycle_a[159] ,rand_second_cycle_a[160] ,rand_second_cycle_a[161] ,rand_second_cycle_a[162] ,rand_second_cycle_a[163] ,rand_second_cycle_a[164] ,rand_second_cycle_a[165] ,rand_second_cycle_a[166] ,rand_second_cycle_a[167] ,rand_second_cycle_a[168] ,rand_second_cycle_a[169] ,rand_second_cycle_a[170] ,rand_second_cycle_a[171] ,rand_second_cycle_a[172] ,rand_second_cycle_a[173] ,rand_second_cycle_a[174] ,rand_second_cycle_a[175] ,rand_second_cycle_a[176] ,rand_second_cycle_a[177] ,rand_second_cycle_a[178] ,rand_second_cycle_a[179] ,rand_second_cycle_a[180] ,rand_second_cycle_a[181] ,rand_second_cycle_a[182] ,rand_second_cycle_a[183] ,rand_second_cycle_a[184] ,rand_second_cycle_a[185] ,rand_second_cycle_a[186] ,rand_second_cycle_a[187] ,rand_second_cycle_a[188] ,rand_second_cycle_a[189] ,rand_second_cycle_a[190] ,rand_second_cycle_a[191] ,rand_second_cycle_a[192] ,rand_second_cycle_a[193] ,rand_second_cycle_a[194] ,rand_second_cycle_a[195] ,rand_second_cycle_a[196] ,rand_second_cycle_a[197] ,rand_second_cycle_a[198] ,rand_second_cycle_a[199] ,rand_second_cycle_a[200] ,rand_second_cycle_a[201] ,rand_second_cycle_a[202] ,rand_second_cycle_a[203] ,rand_second_cycle_a[204] ,rand_second_cycle_a[205] ,rand_second_cycle_a[206] ,rand_second_cycle_a[207] ,rand_second_cycle_a[208] ,rand_second_cycle_a[209] ,rand_second_cycle_a[210] ,rand_second_cycle_a[211] ,rand_second_cycle_a[212] ,rand_second_cycle_a[213] ,rand_second_cycle_a[214] ,rand_second_cycle_a[215] ,rand_second_cycle_a[216] ,rand_second_cycle_a[217] ,rand_second_cycle_a[218] ,rand_second_cycle_a[219] ,rand_second_cycle_a[220] ,rand_second_cycle_a[221] ,rand_second_cycle_a[222] ,rand_second_cycle_a[223] ,rand_second_cycle_a[224] ,rand_second_cycle_a[225] ,rand_second_cycle_a[226] ,rand_second_cycle_a[227] ,rand_second_cycle_a[228] ,rand_second_cycle_a[229] ,rand_second_cycle_a[230] ,rand_second_cycle_a[231] ,rand_second_cycle_a[232] ,rand_second_cycle_a[233] ,rand_second_cycle_a[234] ,rand_second_cycle_a[235] ,rand_second_cycle_a[236] ,rand_second_cycle_a[237] ,rand_second_cycle_a[238] ,rand_second_cycle_a[239] ,rand_second_cycle_a[240] ,rand_second_cycle_a[241] ,rand_second_cycle_a[242] ,rand_second_cycle_a[243] ,rand_second_cycle_a[244] ,rand_second_cycle_a[245] ,rand_second_cycle_a[246] ,rand_second_cycle_a[247] ,rand_second_cycle_a[248] ,rand_second_cycle_a[249] ,rand_second_cycle_a[250] ,rand_second_cycle_a[251] ,rand_second_cycle_a[252] ,rand_second_cycle_a[253] ,rand_second_cycle_a[254] ,
    rand_second_cycle_b[1] ,rand_second_cycle_b[2] ,rand_second_cycle_b[3] ,rand_second_cycle_b[4] ,rand_second_cycle_b[5] ,rand_second_cycle_b[6] ,rand_second_cycle_b[7] ,rand_second_cycle_b[8] ,rand_second_cycle_b[9] ,rand_second_cycle_b[10] ,rand_second_cycle_b[11] ,rand_second_cycle_b[12] ,rand_second_cycle_b[13] ,rand_second_cycle_b[14] ,rand_second_cycle_b[15] ,rand_second_cycle_b[16] ,rand_second_cycle_b[17] ,rand_second_cycle_b[18] ,rand_second_cycle_b[19] ,rand_second_cycle_b[20] ,rand_second_cycle_b[21] ,rand_second_cycle_b[22] ,rand_second_cycle_b[23] ,rand_second_cycle_b[24] ,rand_second_cycle_b[25] ,rand_second_cycle_b[26] ,rand_second_cycle_b[27] ,rand_second_cycle_b[28] ,rand_second_cycle_b[29] ,rand_second_cycle_b[30] ,rand_second_cycle_b[31] ,rand_second_cycle_b[32] ,rand_second_cycle_b[33] ,rand_second_cycle_b[34] ,rand_second_cycle_b[35] ,rand_second_cycle_b[36] ,rand_second_cycle_b[37] ,rand_second_cycle_b[38] ,rand_second_cycle_b[39] ,rand_second_cycle_b[40] ,rand_second_cycle_b[41] ,rand_second_cycle_b[42] ,rand_second_cycle_b[43] ,rand_second_cycle_b[44] ,rand_second_cycle_b[45] ,rand_second_cycle_b[46] ,rand_second_cycle_b[47] ,rand_second_cycle_b[48] ,rand_second_cycle_b[49] ,rand_second_cycle_b[50] ,rand_second_cycle_b[51] ,rand_second_cycle_b[52] ,rand_second_cycle_b[53] ,rand_second_cycle_b[54] ,rand_second_cycle_b[55] ,rand_second_cycle_b[56] ,rand_second_cycle_b[57] ,rand_second_cycle_b[58] ,rand_second_cycle_b[59] ,rand_second_cycle_b[60] ,rand_second_cycle_b[61] ,rand_second_cycle_b[62] ,rand_second_cycle_b[63] ,rand_second_cycle_b[64] ,rand_second_cycle_b[65] ,rand_second_cycle_b[66] ,rand_second_cycle_b[67] ,rand_second_cycle_b[68] ,rand_second_cycle_b[69] ,rand_second_cycle_b[70] ,rand_second_cycle_b[71] ,rand_second_cycle_b[72] ,rand_second_cycle_b[73] ,rand_second_cycle_b[74] ,rand_second_cycle_b[75] ,rand_second_cycle_b[76] ,rand_second_cycle_b[77] ,rand_second_cycle_b[78] ,rand_second_cycle_b[79] ,rand_second_cycle_b[80] ,rand_second_cycle_b[81] ,rand_second_cycle_b[82] ,rand_second_cycle_b[83] ,rand_second_cycle_b[84] ,rand_second_cycle_b[85] ,rand_second_cycle_b[86] ,rand_second_cycle_b[87] ,rand_second_cycle_b[88] ,rand_second_cycle_b[89] ,rand_second_cycle_b[90] ,rand_second_cycle_b[91] ,rand_second_cycle_b[92] ,rand_second_cycle_b[93] ,rand_second_cycle_b[94] ,rand_second_cycle_b[95] ,rand_second_cycle_b[96] ,rand_second_cycle_b[97] ,rand_second_cycle_b[98] ,rand_second_cycle_b[99] ,rand_second_cycle_b[100] ,rand_second_cycle_b[101] ,rand_second_cycle_b[102] ,rand_second_cycle_b[103] ,rand_second_cycle_b[104] ,rand_second_cycle_b[105] ,rand_second_cycle_b[106] ,rand_second_cycle_b[107] ,rand_second_cycle_b[108] ,rand_second_cycle_b[109] ,rand_second_cycle_b[110] ,rand_second_cycle_b[111] ,rand_second_cycle_b[112] ,rand_second_cycle_b[113] ,rand_second_cycle_b[114] ,rand_second_cycle_b[115] ,rand_second_cycle_b[116] ,rand_second_cycle_b[117] ,rand_second_cycle_b[118] ,rand_second_cycle_b[119] ,rand_second_cycle_b[120] ,rand_second_cycle_b[121] ,rand_second_cycle_b[122] ,rand_second_cycle_b[123] ,rand_second_cycle_b[124] ,rand_second_cycle_b[125] ,rand_second_cycle_b[126] ,rand_second_cycle_b[127] ,rand_second_cycle_b[128] ,rand_second_cycle_b[129] ,rand_second_cycle_b[130] ,rand_second_cycle_b[131] ,rand_second_cycle_b[132] ,rand_second_cycle_b[133] ,rand_second_cycle_b[134] ,rand_second_cycle_b[135] ,rand_second_cycle_b[136] ,rand_second_cycle_b[137] ,rand_second_cycle_b[138] ,rand_second_cycle_b[139] ,rand_second_cycle_b[140] ,rand_second_cycle_b[141] ,rand_second_cycle_b[142] ,rand_second_cycle_b[143] ,rand_second_cycle_b[144] ,rand_second_cycle_b[145] ,rand_second_cycle_b[146] ,rand_second_cycle_b[147] ,rand_second_cycle_b[148] ,rand_second_cycle_b[149] ,rand_second_cycle_b[150] ,rand_second_cycle_b[151] ,rand_second_cycle_b[152] ,rand_second_cycle_b[153] ,rand_second_cycle_b[154] ,rand_second_cycle_b[155] ,rand_second_cycle_b[156] ,rand_second_cycle_b[157] ,rand_second_cycle_b[158] ,rand_second_cycle_b[159] ,rand_second_cycle_b[160] ,rand_second_cycle_b[161] ,rand_second_cycle_b[162] ,rand_second_cycle_b[163] ,rand_second_cycle_b[164] ,rand_second_cycle_b[165] ,rand_second_cycle_b[166] ,rand_second_cycle_b[167] ,rand_second_cycle_b[168] ,rand_second_cycle_b[169] ,rand_second_cycle_b[170] ,rand_second_cycle_b[171] ,rand_second_cycle_b[172] ,rand_second_cycle_b[173] ,rand_second_cycle_b[174] ,rand_second_cycle_b[175] ,rand_second_cycle_b[176] ,rand_second_cycle_b[177] ,rand_second_cycle_b[178] ,rand_second_cycle_b[179] ,rand_second_cycle_b[180] ,rand_second_cycle_b[181] ,rand_second_cycle_b[182] ,rand_second_cycle_b[183] ,rand_second_cycle_b[184] ,rand_second_cycle_b[185] ,rand_second_cycle_b[186] ,rand_second_cycle_b[187] ,rand_second_cycle_b[188] ,rand_second_cycle_b[189] ,rand_second_cycle_b[190] ,rand_second_cycle_b[191] ,rand_second_cycle_b[192] ,rand_second_cycle_b[193] ,rand_second_cycle_b[194] ,rand_second_cycle_b[195] ,rand_second_cycle_b[196] ,rand_second_cycle_b[197] ,rand_second_cycle_b[198] ,rand_second_cycle_b[199] ,rand_second_cycle_b[200] ,rand_second_cycle_b[201] ,rand_second_cycle_b[202] ,rand_second_cycle_b[203] ,rand_second_cycle_b[204] ,rand_second_cycle_b[205] ,rand_second_cycle_b[206] ,rand_second_cycle_b[207] ,rand_second_cycle_b[208] ,rand_second_cycle_b[209] ,rand_second_cycle_b[210] ,rand_second_cycle_b[211] ,rand_second_cycle_b[212] ,rand_second_cycle_b[213] ,rand_second_cycle_b[214] ,rand_second_cycle_b[215] ,rand_second_cycle_b[216] ,rand_second_cycle_b[217] ,rand_second_cycle_b[218] ,rand_second_cycle_b[219] ,rand_second_cycle_b[220] ,rand_second_cycle_b[221] ,rand_second_cycle_b[222] ,rand_second_cycle_b[223] ,rand_second_cycle_b[224] ,rand_second_cycle_b[225] ,rand_second_cycle_b[226] ,rand_second_cycle_b[227] ,rand_second_cycle_b[228] ,rand_second_cycle_b[229] ,rand_second_cycle_b[230] ,rand_second_cycle_b[231] ,rand_second_cycle_b[232] ,rand_second_cycle_b[233] ,rand_second_cycle_b[234] ,rand_second_cycle_b[235] ,rand_second_cycle_b[236] ,rand_second_cycle_b[237] ,rand_second_cycle_b[238] ,rand_second_cycle_b[239] ,rand_second_cycle_b[240] ,rand_second_cycle_b[241] ,rand_second_cycle_b[242] ,rand_second_cycle_b[243] ,rand_second_cycle_b[244] ,rand_second_cycle_b[245] ,rand_second_cycle_b[246] ,rand_second_cycle_b[247] ,rand_second_cycle_b[248] ,rand_second_cycle_b[249] ,rand_second_cycle_b[250] ,rand_second_cycle_b[251] ,rand_second_cycle_b[252] ,rand_second_cycle_b[253] ,rand_second_cycle_b[254] ,
    x0_subscript1_share3_wire, x1_subscript1_share3_wire, x2_subscript1_share3_wire, x3_subscript1_share3_wire, x4_subscript1_share3_wire, x5_subscript1_share3_wire, x6_subscript1_share3_wire, x7_subscript1_share3_wire , x0x1_subscript1_share3_wire , x0x2_subscript1_share3_wire , x0x3_subscript1_share3_wire , x0x4_subscript1_share3_wire , x0x5_subscript1_share3_wire , x0x6_subscript1_share3_wire , x0x7_subscript1_share3_wire , x1x2_subscript1_share3_wire , x1x3_subscript1_share3_wire , x1x4_subscript1_share3_wire , x1x5_subscript1_share3_wire , x1x6_subscript1_share3_wire , x1x7_subscript1_share3_wire , x2x3_subscript1_share3_wire , x2x4_subscript1_share3_wire , x2x5_subscript1_share3_wire , x2x6_subscript1_share3_wire , x2x7_subscript1_share3_wire , x3x4_subscript1_share3_wire , x3x5_subscript1_share3_wire , x3x6_subscript1_share3_wire , x3x7_subscript1_share3_wire , x4x5_subscript1_share3_wire , x4x6_subscript1_share3_wire , x4x7_subscript1_share3_wire , x5x6_subscript1_share3_wire , x5x7_subscript1_share3_wire , x6x7_subscript1_share3_wire , x0x1x2_subscript1_share3_wire , x0x1x3_subscript1_share3_wire , x0x1x4_subscript1_share3_wire , x0x1x5_subscript1_share3_wire , x0x1x6_subscript1_share3_wire , x0x1x7_subscript1_share3_wire , x0x2x3_subscript1_share3_wire , x0x2x4_subscript1_share3_wire , x0x2x5_subscript1_share3_wire , x0x2x6_subscript1_share3_wire , x0x2x7_subscript1_share3_wire , x0x3x4_subscript1_share3_wire , x0x3x5_subscript1_share3_wire , x0x3x6_subscript1_share3_wire , x0x3x7_subscript1_share3_wire , x0x4x5_subscript1_share3_wire , x0x4x6_subscript1_share3_wire , x0x4x7_subscript1_share3_wire , x0x5x6_subscript1_share3_wire , x0x5x7_subscript1_share3_wire , x0x6x7_subscript1_share3_wire , x1x2x3_subscript1_share3_wire , x1x2x4_subscript1_share3_wire , x1x2x5_subscript1_share3_wire , x1x2x6_subscript1_share3_wire , x1x2x7_subscript1_share3_wire , x1x3x4_subscript1_share3_wire , x1x3x5_subscript1_share3_wire , x1x3x6_subscript1_share3_wire , x1x3x7_subscript1_share3_wire , x1x4x5_subscript1_share3_wire , x1x4x6_subscript1_share3_wire , x1x4x7_subscript1_share3_wire , x1x5x6_subscript1_share3_wire , x1x5x7_subscript1_share3_wire , x1x6x7_subscript1_share3_wire , x2x3x4_subscript1_share3_wire , x2x3x5_subscript1_share3_wire , x2x3x6_subscript1_share3_wire , x2x3x7_subscript1_share3_wire , x2x4x5_subscript1_share3_wire , x2x4x6_subscript1_share3_wire , x2x4x7_subscript1_share3_wire , x2x5x6_subscript1_share3_wire , x2x5x7_subscript1_share3_wire , x2x6x7_subscript1_share3_wire , x3x4x5_subscript1_share3_wire , x3x4x6_subscript1_share3_wire , x3x4x7_subscript1_share3_wire , x3x5x6_subscript1_share3_wire , x3x5x7_subscript1_share3_wire , x3x6x7_subscript1_share3_wire , x4x5x6_subscript1_share3_wire , x4x5x7_subscript1_share3_wire , x4x6x7_subscript1_share3_wire , x5x6x7_subscript1_share3_wire , x0x1x2x3_subscript1_share3_wire , x0x1x2x4_subscript1_share3_wire , x0x1x2x5_subscript1_share3_wire , x0x1x2x6_subscript1_share3_wire , x0x1x2x7_subscript1_share3_wire , x0x1x3x4_subscript1_share3_wire , x0x1x3x5_subscript1_share3_wire , x0x1x3x6_subscript1_share3_wire , x0x1x3x7_subscript1_share3_wire , x0x1x4x5_subscript1_share3_wire , x0x1x4x6_subscript1_share3_wire , x0x1x4x7_subscript1_share3_wire , x0x1x5x6_subscript1_share3_wire , x0x1x5x7_subscript1_share3_wire , x0x1x6x7_subscript1_share3_wire , x0x2x3x4_subscript1_share3_wire , x0x2x3x5_subscript1_share3_wire , x0x2x3x6_subscript1_share3_wire , x0x2x3x7_subscript1_share3_wire , x0x2x4x5_subscript1_share3_wire , x0x2x4x6_subscript1_share3_wire , x0x2x4x7_subscript1_share3_wire , x0x2x5x6_subscript1_share3_wire , x0x2x5x7_subscript1_share3_wire , x0x2x6x7_subscript1_share3_wire , x0x3x4x5_subscript1_share3_wire , x0x3x4x6_subscript1_share3_wire , x0x3x4x7_subscript1_share3_wire , x0x3x5x6_subscript1_share3_wire , x0x3x5x7_subscript1_share3_wire , x0x3x6x7_subscript1_share3_wire , x0x4x5x6_subscript1_share3_wire , x0x4x5x7_subscript1_share3_wire , x0x4x6x7_subscript1_share3_wire , x0x5x6x7_subscript1_share3_wire , x1x2x3x4_subscript1_share3_wire , x1x2x3x5_subscript1_share3_wire , x1x2x3x6_subscript1_share3_wire , x1x2x3x7_subscript1_share3_wire , x1x2x4x5_subscript1_share3_wire , x1x2x4x6_subscript1_share3_wire , x1x2x4x7_subscript1_share3_wire , x1x2x5x6_subscript1_share3_wire , x1x2x5x7_subscript1_share3_wire , x1x2x6x7_subscript1_share3_wire , x1x3x4x5_subscript1_share3_wire , x1x3x4x6_subscript1_share3_wire , x1x3x4x7_subscript1_share3_wire , x1x3x5x6_subscript1_share3_wire , x1x3x5x7_subscript1_share3_wire , x1x3x6x7_subscript1_share3_wire , x1x4x5x6_subscript1_share3_wire , x1x4x5x7_subscript1_share3_wire , x1x4x6x7_subscript1_share3_wire , x1x5x6x7_subscript1_share3_wire , x2x3x4x5_subscript1_share3_wire , x2x3x4x6_subscript1_share3_wire , x2x3x4x7_subscript1_share3_wire , x2x3x5x6_subscript1_share3_wire , x2x3x5x7_subscript1_share3_wire , x2x3x6x7_subscript1_share3_wire , x2x4x5x6_subscript1_share3_wire , x2x4x5x7_subscript1_share3_wire , x2x4x6x7_subscript1_share3_wire , x2x5x6x7_subscript1_share3_wire , x3x4x5x6_subscript1_share3_wire , x3x4x5x7_subscript1_share3_wire , x3x4x6x7_subscript1_share3_wire , x3x5x6x7_subscript1_share3_wire , x4x5x6x7_subscript1_share3_wire , x0x1x2x3x4_subscript1_share3_wire , x0x1x2x3x5_subscript1_share3_wire , x0x1x2x3x6_subscript1_share3_wire , x0x1x2x3x7_subscript1_share3_wire , x0x1x2x4x5_subscript1_share3_wire , x0x1x2x4x6_subscript1_share3_wire , x0x1x2x4x7_subscript1_share3_wire , x0x1x2x5x6_subscript1_share3_wire , x0x1x2x5x7_subscript1_share3_wire , x0x1x2x6x7_subscript1_share3_wire , x0x1x3x4x5_subscript1_share3_wire , x0x1x3x4x6_subscript1_share3_wire , x0x1x3x4x7_subscript1_share3_wire , x0x1x3x5x6_subscript1_share3_wire , x0x1x3x5x7_subscript1_share3_wire , x0x1x3x6x7_subscript1_share3_wire , x0x1x4x5x6_subscript1_share3_wire , x0x1x4x5x7_subscript1_share3_wire , x0x1x4x6x7_subscript1_share3_wire , x0x1x5x6x7_subscript1_share3_wire , x0x2x3x4x5_subscript1_share3_wire , x0x2x3x4x6_subscript1_share3_wire , x0x2x3x4x7_subscript1_share3_wire , x0x2x3x5x6_subscript1_share3_wire , x0x2x3x5x7_subscript1_share3_wire , x0x2x3x6x7_subscript1_share3_wire , x0x2x4x5x6_subscript1_share3_wire , x0x2x4x5x7_subscript1_share3_wire , x0x2x4x6x7_subscript1_share3_wire , x0x2x5x6x7_subscript1_share3_wire , x0x3x4x5x6_subscript1_share3_wire , x0x3x4x5x7_subscript1_share3_wire , x0x3x4x6x7_subscript1_share3_wire , x0x3x5x6x7_subscript1_share3_wire , x0x4x5x6x7_subscript1_share3_wire , x1x2x3x4x5_subscript1_share3_wire , x1x2x3x4x6_subscript1_share3_wire , x1x2x3x4x7_subscript1_share3_wire , x1x2x3x5x6_subscript1_share3_wire , x1x2x3x5x7_subscript1_share3_wire , x1x2x3x6x7_subscript1_share3_wire , x1x2x4x5x6_subscript1_share3_wire , x1x2x4x5x7_subscript1_share3_wire , x1x2x4x6x7_subscript1_share3_wire , x1x2x5x6x7_subscript1_share3_wire , x1x3x4x5x6_subscript1_share3_wire , x1x3x4x5x7_subscript1_share3_wire , x1x3x4x6x7_subscript1_share3_wire , x1x3x5x6x7_subscript1_share3_wire , x1x4x5x6x7_subscript1_share3_wire , x2x3x4x5x6_subscript1_share3_wire , x2x3x4x5x7_subscript1_share3_wire , x2x3x4x6x7_subscript1_share3_wire , x2x3x5x6x7_subscript1_share3_wire , x2x4x5x6x7_subscript1_share3_wire , x3x4x5x6x7_subscript1_share3_wire , x0x1x2x3x4x5_subscript1_share3_wire , x0x1x2x3x4x6_subscript1_share3_wire , x0x1x2x3x4x7_subscript1_share3_wire , x0x1x2x3x5x6_subscript1_share3_wire , x0x1x2x3x5x7_subscript1_share3_wire , x0x1x2x3x6x7_subscript1_share3_wire , x0x1x2x4x5x6_subscript1_share3_wire , x0x1x2x4x5x7_subscript1_share3_wire , x0x1x2x4x6x7_subscript1_share3_wire , x0x1x2x5x6x7_subscript1_share3_wire , x0x1x3x4x5x6_subscript1_share3_wire , x0x1x3x4x5x7_subscript1_share3_wire , x0x1x3x4x6x7_subscript1_share3_wire , x0x1x3x5x6x7_subscript1_share3_wire , x0x1x4x5x6x7_subscript1_share3_wire , x0x2x3x4x5x6_subscript1_share3_wire , x0x2x3x4x5x7_subscript1_share3_wire , x0x2x3x4x6x7_subscript1_share3_wire , x0x2x3x5x6x7_subscript1_share3_wire , x0x2x4x5x6x7_subscript1_share3_wire , x0x3x4x5x6x7_subscript1_share3_wire , x1x2x3x4x5x6_subscript1_share3_wire , x1x2x3x4x5x7_subscript1_share3_wire , x1x2x3x4x6x7_subscript1_share3_wire , x1x2x3x5x6x7_subscript1_share3_wire , x1x2x4x5x6x7_subscript1_share3_wire , x1x3x4x5x6x7_subscript1_share3_wire , x2x3x4x5x6x7_subscript1_share3_wire , x0x1x2x3x4x5x6_subscript1_share3_wire , x0x1x2x3x4x5x7_subscript1_share3_wire , x0x1x2x3x4x6x7_subscript1_share3_wire , x0x1x2x3x5x6x7_subscript1_share3_wire , x0x1x2x4x5x6x7_subscript1_share3_wire , x0x1x3x4x5x6x7_subscript1_share3_wire , x0x2x3x4x5x6x7_subscript1_share3_wire , x1x2x3x4x5x6x7_subscript1_share3_wire 
);

// Register stage 

register_array_AES_oneshare second_cycle_share1_reg (
    clk,
    x0_subscript1_share1_wire, x1_subscript1_share1_wire, x2_subscript1_share1_wire, x3_subscript1_share1_wire, x4_subscript1_share1_wire, x5_subscript1_share1_wire, x6_subscript1_share1_wire, x7_subscript1_share1_wire , x0x1_subscript1_share1_wire , x0x2_subscript1_share1_wire , x0x3_subscript1_share1_wire , x0x4_subscript1_share1_wire , x0x5_subscript1_share1_wire , x0x6_subscript1_share1_wire , x0x7_subscript1_share1_wire , x1x2_subscript1_share1_wire , x1x3_subscript1_share1_wire , x1x4_subscript1_share1_wire , x1x5_subscript1_share1_wire , x1x6_subscript1_share1_wire , x1x7_subscript1_share1_wire , x2x3_subscript1_share1_wire , x2x4_subscript1_share1_wire , x2x5_subscript1_share1_wire , x2x6_subscript1_share1_wire , x2x7_subscript1_share1_wire , x3x4_subscript1_share1_wire , x3x5_subscript1_share1_wire , x3x6_subscript1_share1_wire , x3x7_subscript1_share1_wire , x4x5_subscript1_share1_wire , x4x6_subscript1_share1_wire , x4x7_subscript1_share1_wire , x5x6_subscript1_share1_wire , x5x7_subscript1_share1_wire , x6x7_subscript1_share1_wire , x0x1x2_subscript1_share1_wire , x0x1x3_subscript1_share1_wire , x0x1x4_subscript1_share1_wire , x0x1x5_subscript1_share1_wire , x0x1x6_subscript1_share1_wire , x0x1x7_subscript1_share1_wire , x0x2x3_subscript1_share1_wire , x0x2x4_subscript1_share1_wire , x0x2x5_subscript1_share1_wire , x0x2x6_subscript1_share1_wire , x0x2x7_subscript1_share1_wire , x0x3x4_subscript1_share1_wire , x0x3x5_subscript1_share1_wire , x0x3x6_subscript1_share1_wire , x0x3x7_subscript1_share1_wire , x0x4x5_subscript1_share1_wire , x0x4x6_subscript1_share1_wire , x0x4x7_subscript1_share1_wire , x0x5x6_subscript1_share1_wire , x0x5x7_subscript1_share1_wire , x0x6x7_subscript1_share1_wire , x1x2x3_subscript1_share1_wire , x1x2x4_subscript1_share1_wire , x1x2x5_subscript1_share1_wire , x1x2x6_subscript1_share1_wire , x1x2x7_subscript1_share1_wire , x1x3x4_subscript1_share1_wire , x1x3x5_subscript1_share1_wire , x1x3x6_subscript1_share1_wire , x1x3x7_subscript1_share1_wire , x1x4x5_subscript1_share1_wire , x1x4x6_subscript1_share1_wire , x1x4x7_subscript1_share1_wire , x1x5x6_subscript1_share1_wire , x1x5x7_subscript1_share1_wire , x1x6x7_subscript1_share1_wire , x2x3x4_subscript1_share1_wire , x2x3x5_subscript1_share1_wire , x2x3x6_subscript1_share1_wire , x2x3x7_subscript1_share1_wire , x2x4x5_subscript1_share1_wire , x2x4x6_subscript1_share1_wire , x2x4x7_subscript1_share1_wire , x2x5x6_subscript1_share1_wire , x2x5x7_subscript1_share1_wire , x2x6x7_subscript1_share1_wire , x3x4x5_subscript1_share1_wire , x3x4x6_subscript1_share1_wire , x3x4x7_subscript1_share1_wire , x3x5x6_subscript1_share1_wire , x3x5x7_subscript1_share1_wire , x3x6x7_subscript1_share1_wire , x4x5x6_subscript1_share1_wire , x4x5x7_subscript1_share1_wire , x4x6x7_subscript1_share1_wire , x5x6x7_subscript1_share1_wire , x0x1x2x3_subscript1_share1_wire , x0x1x2x4_subscript1_share1_wire , x0x1x2x5_subscript1_share1_wire , x0x1x2x6_subscript1_share1_wire , x0x1x2x7_subscript1_share1_wire , x0x1x3x4_subscript1_share1_wire , x0x1x3x5_subscript1_share1_wire , x0x1x3x6_subscript1_share1_wire , x0x1x3x7_subscript1_share1_wire , x0x1x4x5_subscript1_share1_wire , x0x1x4x6_subscript1_share1_wire , x0x1x4x7_subscript1_share1_wire , x0x1x5x6_subscript1_share1_wire , x0x1x5x7_subscript1_share1_wire , x0x1x6x7_subscript1_share1_wire , x0x2x3x4_subscript1_share1_wire , x0x2x3x5_subscript1_share1_wire , x0x2x3x6_subscript1_share1_wire , x0x2x3x7_subscript1_share1_wire , x0x2x4x5_subscript1_share1_wire , x0x2x4x6_subscript1_share1_wire , x0x2x4x7_subscript1_share1_wire , x0x2x5x6_subscript1_share1_wire , x0x2x5x7_subscript1_share1_wire , x0x2x6x7_subscript1_share1_wire , x0x3x4x5_subscript1_share1_wire , x0x3x4x6_subscript1_share1_wire , x0x3x4x7_subscript1_share1_wire , x0x3x5x6_subscript1_share1_wire , x0x3x5x7_subscript1_share1_wire , x0x3x6x7_subscript1_share1_wire , x0x4x5x6_subscript1_share1_wire , x0x4x5x7_subscript1_share1_wire , x0x4x6x7_subscript1_share1_wire , x0x5x6x7_subscript1_share1_wire , x1x2x3x4_subscript1_share1_wire , x1x2x3x5_subscript1_share1_wire , x1x2x3x6_subscript1_share1_wire , x1x2x3x7_subscript1_share1_wire , x1x2x4x5_subscript1_share1_wire , x1x2x4x6_subscript1_share1_wire , x1x2x4x7_subscript1_share1_wire , x1x2x5x6_subscript1_share1_wire , x1x2x5x7_subscript1_share1_wire , x1x2x6x7_subscript1_share1_wire , x1x3x4x5_subscript1_share1_wire , x1x3x4x6_subscript1_share1_wire , x1x3x4x7_subscript1_share1_wire , x1x3x5x6_subscript1_share1_wire , x1x3x5x7_subscript1_share1_wire , x1x3x6x7_subscript1_share1_wire , x1x4x5x6_subscript1_share1_wire , x1x4x5x7_subscript1_share1_wire , x1x4x6x7_subscript1_share1_wire , x1x5x6x7_subscript1_share1_wire , x2x3x4x5_subscript1_share1_wire , x2x3x4x6_subscript1_share1_wire , x2x3x4x7_subscript1_share1_wire , x2x3x5x6_subscript1_share1_wire , x2x3x5x7_subscript1_share1_wire , x2x3x6x7_subscript1_share1_wire , x2x4x5x6_subscript1_share1_wire , x2x4x5x7_subscript1_share1_wire , x2x4x6x7_subscript1_share1_wire , x2x5x6x7_subscript1_share1_wire , x3x4x5x6_subscript1_share1_wire , x3x4x5x7_subscript1_share1_wire , x3x4x6x7_subscript1_share1_wire , x3x5x6x7_subscript1_share1_wire , x4x5x6x7_subscript1_share1_wire , x0x1x2x3x4_subscript1_share1_wire , x0x1x2x3x5_subscript1_share1_wire , x0x1x2x3x6_subscript1_share1_wire , x0x1x2x3x7_subscript1_share1_wire , x0x1x2x4x5_subscript1_share1_wire , x0x1x2x4x6_subscript1_share1_wire , x0x1x2x4x7_subscript1_share1_wire , x0x1x2x5x6_subscript1_share1_wire , x0x1x2x5x7_subscript1_share1_wire , x0x1x2x6x7_subscript1_share1_wire , x0x1x3x4x5_subscript1_share1_wire , x0x1x3x4x6_subscript1_share1_wire , x0x1x3x4x7_subscript1_share1_wire , x0x1x3x5x6_subscript1_share1_wire , x0x1x3x5x7_subscript1_share1_wire , x0x1x3x6x7_subscript1_share1_wire , x0x1x4x5x6_subscript1_share1_wire , x0x1x4x5x7_subscript1_share1_wire , x0x1x4x6x7_subscript1_share1_wire , x0x1x5x6x7_subscript1_share1_wire , x0x2x3x4x5_subscript1_share1_wire , x0x2x3x4x6_subscript1_share1_wire , x0x2x3x4x7_subscript1_share1_wire , x0x2x3x5x6_subscript1_share1_wire , x0x2x3x5x7_subscript1_share1_wire , x0x2x3x6x7_subscript1_share1_wire , x0x2x4x5x6_subscript1_share1_wire , x0x2x4x5x7_subscript1_share1_wire , x0x2x4x6x7_subscript1_share1_wire , x0x2x5x6x7_subscript1_share1_wire , x0x3x4x5x6_subscript1_share1_wire , x0x3x4x5x7_subscript1_share1_wire , x0x3x4x6x7_subscript1_share1_wire , x0x3x5x6x7_subscript1_share1_wire , x0x4x5x6x7_subscript1_share1_wire , x1x2x3x4x5_subscript1_share1_wire , x1x2x3x4x6_subscript1_share1_wire , x1x2x3x4x7_subscript1_share1_wire , x1x2x3x5x6_subscript1_share1_wire , x1x2x3x5x7_subscript1_share1_wire , x1x2x3x6x7_subscript1_share1_wire , x1x2x4x5x6_subscript1_share1_wire , x1x2x4x5x7_subscript1_share1_wire , x1x2x4x6x7_subscript1_share1_wire , x1x2x5x6x7_subscript1_share1_wire , x1x3x4x5x6_subscript1_share1_wire , x1x3x4x5x7_subscript1_share1_wire , x1x3x4x6x7_subscript1_share1_wire , x1x3x5x6x7_subscript1_share1_wire , x1x4x5x6x7_subscript1_share1_wire , x2x3x4x5x6_subscript1_share1_wire , x2x3x4x5x7_subscript1_share1_wire , x2x3x4x6x7_subscript1_share1_wire , x2x3x5x6x7_subscript1_share1_wire , x2x4x5x6x7_subscript1_share1_wire , x3x4x5x6x7_subscript1_share1_wire , x0x1x2x3x4x5_subscript1_share1_wire , x0x1x2x3x4x6_subscript1_share1_wire , x0x1x2x3x4x7_subscript1_share1_wire , x0x1x2x3x5x6_subscript1_share1_wire , x0x1x2x3x5x7_subscript1_share1_wire , x0x1x2x3x6x7_subscript1_share1_wire , x0x1x2x4x5x6_subscript1_share1_wire , x0x1x2x4x5x7_subscript1_share1_wire , x0x1x2x4x6x7_subscript1_share1_wire , x0x1x2x5x6x7_subscript1_share1_wire , x0x1x3x4x5x6_subscript1_share1_wire , x0x1x3x4x5x7_subscript1_share1_wire , x0x1x3x4x6x7_subscript1_share1_wire , x0x1x3x5x6x7_subscript1_share1_wire , x0x1x4x5x6x7_subscript1_share1_wire , x0x2x3x4x5x6_subscript1_share1_wire , x0x2x3x4x5x7_subscript1_share1_wire , x0x2x3x4x6x7_subscript1_share1_wire , x0x2x3x5x6x7_subscript1_share1_wire , x0x2x4x5x6x7_subscript1_share1_wire , x0x3x4x5x6x7_subscript1_share1_wire , x1x2x3x4x5x6_subscript1_share1_wire , x1x2x3x4x5x7_subscript1_share1_wire , x1x2x3x4x6x7_subscript1_share1_wire , x1x2x3x5x6x7_subscript1_share1_wire , x1x2x4x5x6x7_subscript1_share1_wire , x1x3x4x5x6x7_subscript1_share1_wire , x2x3x4x5x6x7_subscript1_share1_wire , x0x1x2x3x4x5x6_subscript1_share1_wire , x0x1x2x3x4x5x7_subscript1_share1_wire , x0x1x2x3x4x6x7_subscript1_share1_wire , x0x1x2x3x5x6x7_subscript1_share1_wire , x0x1x2x4x5x6x7_subscript1_share1_wire , x0x1x3x4x5x6x7_subscript1_share1_wire , x0x2x3x4x5x6x7_subscript1_share1_wire , x1x2x3x4x5x6x7_subscript1_share1_wire ,
    x0_subscript1_share1_reg, x1_subscript1_share1_reg, x2_subscript1_share1_reg, x3_subscript1_share1_reg, x4_subscript1_share1_reg, x5_subscript1_share1_reg, x6_subscript1_share1_reg, x7_subscript1_share1_reg , x0x1_subscript1_share1_reg , x0x2_subscript1_share1_reg , x0x3_subscript1_share1_reg , x0x4_subscript1_share1_reg , x0x5_subscript1_share1_reg , x0x6_subscript1_share1_reg , x0x7_subscript1_share1_reg , x1x2_subscript1_share1_reg , x1x3_subscript1_share1_reg , x1x4_subscript1_share1_reg , x1x5_subscript1_share1_reg , x1x6_subscript1_share1_reg , x1x7_subscript1_share1_reg , x2x3_subscript1_share1_reg , x2x4_subscript1_share1_reg , x2x5_subscript1_share1_reg , x2x6_subscript1_share1_reg , x2x7_subscript1_share1_reg , x3x4_subscript1_share1_reg , x3x5_subscript1_share1_reg , x3x6_subscript1_share1_reg , x3x7_subscript1_share1_reg , x4x5_subscript1_share1_reg , x4x6_subscript1_share1_reg , x4x7_subscript1_share1_reg , x5x6_subscript1_share1_reg , x5x7_subscript1_share1_reg , x6x7_subscript1_share1_reg , x0x1x2_subscript1_share1_reg , x0x1x3_subscript1_share1_reg , x0x1x4_subscript1_share1_reg , x0x1x5_subscript1_share1_reg , x0x1x6_subscript1_share1_reg , x0x1x7_subscript1_share1_reg , x0x2x3_subscript1_share1_reg , x0x2x4_subscript1_share1_reg , x0x2x5_subscript1_share1_reg , x0x2x6_subscript1_share1_reg , x0x2x7_subscript1_share1_reg , x0x3x4_subscript1_share1_reg , x0x3x5_subscript1_share1_reg , x0x3x6_subscript1_share1_reg , x0x3x7_subscript1_share1_reg , x0x4x5_subscript1_share1_reg , x0x4x6_subscript1_share1_reg , x0x4x7_subscript1_share1_reg , x0x5x6_subscript1_share1_reg , x0x5x7_subscript1_share1_reg , x0x6x7_subscript1_share1_reg , x1x2x3_subscript1_share1_reg , x1x2x4_subscript1_share1_reg , x1x2x5_subscript1_share1_reg , x1x2x6_subscript1_share1_reg , x1x2x7_subscript1_share1_reg , x1x3x4_subscript1_share1_reg , x1x3x5_subscript1_share1_reg , x1x3x6_subscript1_share1_reg , x1x3x7_subscript1_share1_reg , x1x4x5_subscript1_share1_reg , x1x4x6_subscript1_share1_reg , x1x4x7_subscript1_share1_reg , x1x5x6_subscript1_share1_reg , x1x5x7_subscript1_share1_reg , x1x6x7_subscript1_share1_reg , x2x3x4_subscript1_share1_reg , x2x3x5_subscript1_share1_reg , x2x3x6_subscript1_share1_reg , x2x3x7_subscript1_share1_reg , x2x4x5_subscript1_share1_reg , x2x4x6_subscript1_share1_reg , x2x4x7_subscript1_share1_reg , x2x5x6_subscript1_share1_reg , x2x5x7_subscript1_share1_reg , x2x6x7_subscript1_share1_reg , x3x4x5_subscript1_share1_reg , x3x4x6_subscript1_share1_reg , x3x4x7_subscript1_share1_reg , x3x5x6_subscript1_share1_reg , x3x5x7_subscript1_share1_reg , x3x6x7_subscript1_share1_reg , x4x5x6_subscript1_share1_reg , x4x5x7_subscript1_share1_reg , x4x6x7_subscript1_share1_reg , x5x6x7_subscript1_share1_reg , x0x1x2x3_subscript1_share1_reg , x0x1x2x4_subscript1_share1_reg , x0x1x2x5_subscript1_share1_reg , x0x1x2x6_subscript1_share1_reg , x0x1x2x7_subscript1_share1_reg , x0x1x3x4_subscript1_share1_reg , x0x1x3x5_subscript1_share1_reg , x0x1x3x6_subscript1_share1_reg , x0x1x3x7_subscript1_share1_reg , x0x1x4x5_subscript1_share1_reg , x0x1x4x6_subscript1_share1_reg , x0x1x4x7_subscript1_share1_reg , x0x1x5x6_subscript1_share1_reg , x0x1x5x7_subscript1_share1_reg , x0x1x6x7_subscript1_share1_reg , x0x2x3x4_subscript1_share1_reg , x0x2x3x5_subscript1_share1_reg , x0x2x3x6_subscript1_share1_reg , x0x2x3x7_subscript1_share1_reg , x0x2x4x5_subscript1_share1_reg , x0x2x4x6_subscript1_share1_reg , x0x2x4x7_subscript1_share1_reg , x0x2x5x6_subscript1_share1_reg , x0x2x5x7_subscript1_share1_reg , x0x2x6x7_subscript1_share1_reg , x0x3x4x5_subscript1_share1_reg , x0x3x4x6_subscript1_share1_reg , x0x3x4x7_subscript1_share1_reg , x0x3x5x6_subscript1_share1_reg , x0x3x5x7_subscript1_share1_reg , x0x3x6x7_subscript1_share1_reg , x0x4x5x6_subscript1_share1_reg , x0x4x5x7_subscript1_share1_reg , x0x4x6x7_subscript1_share1_reg , x0x5x6x7_subscript1_share1_reg , x1x2x3x4_subscript1_share1_reg , x1x2x3x5_subscript1_share1_reg , x1x2x3x6_subscript1_share1_reg , x1x2x3x7_subscript1_share1_reg , x1x2x4x5_subscript1_share1_reg , x1x2x4x6_subscript1_share1_reg , x1x2x4x7_subscript1_share1_reg , x1x2x5x6_subscript1_share1_reg , x1x2x5x7_subscript1_share1_reg , x1x2x6x7_subscript1_share1_reg , x1x3x4x5_subscript1_share1_reg , x1x3x4x6_subscript1_share1_reg , x1x3x4x7_subscript1_share1_reg , x1x3x5x6_subscript1_share1_reg , x1x3x5x7_subscript1_share1_reg , x1x3x6x7_subscript1_share1_reg , x1x4x5x6_subscript1_share1_reg , x1x4x5x7_subscript1_share1_reg , x1x4x6x7_subscript1_share1_reg , x1x5x6x7_subscript1_share1_reg , x2x3x4x5_subscript1_share1_reg , x2x3x4x6_subscript1_share1_reg , x2x3x4x7_subscript1_share1_reg , x2x3x5x6_subscript1_share1_reg , x2x3x5x7_subscript1_share1_reg , x2x3x6x7_subscript1_share1_reg , x2x4x5x6_subscript1_share1_reg , x2x4x5x7_subscript1_share1_reg , x2x4x6x7_subscript1_share1_reg , x2x5x6x7_subscript1_share1_reg , x3x4x5x6_subscript1_share1_reg , x3x4x5x7_subscript1_share1_reg , x3x4x6x7_subscript1_share1_reg , x3x5x6x7_subscript1_share1_reg , x4x5x6x7_subscript1_share1_reg , x0x1x2x3x4_subscript1_share1_reg , x0x1x2x3x5_subscript1_share1_reg , x0x1x2x3x6_subscript1_share1_reg , x0x1x2x3x7_subscript1_share1_reg , x0x1x2x4x5_subscript1_share1_reg , x0x1x2x4x6_subscript1_share1_reg , x0x1x2x4x7_subscript1_share1_reg , x0x1x2x5x6_subscript1_share1_reg , x0x1x2x5x7_subscript1_share1_reg , x0x1x2x6x7_subscript1_share1_reg , x0x1x3x4x5_subscript1_share1_reg , x0x1x3x4x6_subscript1_share1_reg , x0x1x3x4x7_subscript1_share1_reg , x0x1x3x5x6_subscript1_share1_reg , x0x1x3x5x7_subscript1_share1_reg , x0x1x3x6x7_subscript1_share1_reg , x0x1x4x5x6_subscript1_share1_reg , x0x1x4x5x7_subscript1_share1_reg , x0x1x4x6x7_subscript1_share1_reg , x0x1x5x6x7_subscript1_share1_reg , x0x2x3x4x5_subscript1_share1_reg , x0x2x3x4x6_subscript1_share1_reg , x0x2x3x4x7_subscript1_share1_reg , x0x2x3x5x6_subscript1_share1_reg , x0x2x3x5x7_subscript1_share1_reg , x0x2x3x6x7_subscript1_share1_reg , x0x2x4x5x6_subscript1_share1_reg , x0x2x4x5x7_subscript1_share1_reg , x0x2x4x6x7_subscript1_share1_reg , x0x2x5x6x7_subscript1_share1_reg , x0x3x4x5x6_subscript1_share1_reg , x0x3x4x5x7_subscript1_share1_reg , x0x3x4x6x7_subscript1_share1_reg , x0x3x5x6x7_subscript1_share1_reg , x0x4x5x6x7_subscript1_share1_reg , x1x2x3x4x5_subscript1_share1_reg , x1x2x3x4x6_subscript1_share1_reg , x1x2x3x4x7_subscript1_share1_reg , x1x2x3x5x6_subscript1_share1_reg , x1x2x3x5x7_subscript1_share1_reg , x1x2x3x6x7_subscript1_share1_reg , x1x2x4x5x6_subscript1_share1_reg , x1x2x4x5x7_subscript1_share1_reg , x1x2x4x6x7_subscript1_share1_reg , x1x2x5x6x7_subscript1_share1_reg , x1x3x4x5x6_subscript1_share1_reg , x1x3x4x5x7_subscript1_share1_reg , x1x3x4x6x7_subscript1_share1_reg , x1x3x5x6x7_subscript1_share1_reg , x1x4x5x6x7_subscript1_share1_reg , x2x3x4x5x6_subscript1_share1_reg , x2x3x4x5x7_subscript1_share1_reg , x2x3x4x6x7_subscript1_share1_reg , x2x3x5x6x7_subscript1_share1_reg , x2x4x5x6x7_subscript1_share1_reg , x3x4x5x6x7_subscript1_share1_reg , x0x1x2x3x4x5_subscript1_share1_reg , x0x1x2x3x4x6_subscript1_share1_reg , x0x1x2x3x4x7_subscript1_share1_reg , x0x1x2x3x5x6_subscript1_share1_reg , x0x1x2x3x5x7_subscript1_share1_reg , x0x1x2x3x6x7_subscript1_share1_reg , x0x1x2x4x5x6_subscript1_share1_reg , x0x1x2x4x5x7_subscript1_share1_reg , x0x1x2x4x6x7_subscript1_share1_reg , x0x1x2x5x6x7_subscript1_share1_reg , x0x1x3x4x5x6_subscript1_share1_reg , x0x1x3x4x5x7_subscript1_share1_reg , x0x1x3x4x6x7_subscript1_share1_reg , x0x1x3x5x6x7_subscript1_share1_reg , x0x1x4x5x6x7_subscript1_share1_reg , x0x2x3x4x5x6_subscript1_share1_reg , x0x2x3x4x5x7_subscript1_share1_reg , x0x2x3x4x6x7_subscript1_share1_reg , x0x2x3x5x6x7_subscript1_share1_reg , x0x2x4x5x6x7_subscript1_share1_reg , x0x3x4x5x6x7_subscript1_share1_reg , x1x2x3x4x5x6_subscript1_share1_reg , x1x2x3x4x5x7_subscript1_share1_reg , x1x2x3x4x6x7_subscript1_share1_reg , x1x2x3x5x6x7_subscript1_share1_reg , x1x2x4x5x6x7_subscript1_share1_reg , x1x3x4x5x6x7_subscript1_share1_reg , x2x3x4x5x6x7_subscript1_share1_reg , x0x1x2x3x4x5x6_subscript1_share1_reg , x0x1x2x3x4x5x7_subscript1_share1_reg , x0x1x2x3x4x6x7_subscript1_share1_reg , x0x1x2x3x5x6x7_subscript1_share1_reg , x0x1x2x4x5x6x7_subscript1_share1_reg , x0x1x3x4x5x6x7_subscript1_share1_reg , x0x2x3x4x5x6x7_subscript1_share1_reg , x1x2x3x4x5x6x7_subscript1_share1_reg 
);
register_array_AES_oneshare second_cycle_share2_reg (
    clk,
    x0_subscript1_share2_wire, x1_subscript1_share2_wire, x2_subscript1_share2_wire, x3_subscript1_share2_wire, x4_subscript1_share2_wire, x5_subscript1_share2_wire, x6_subscript1_share2_wire, x7_subscript1_share2_wire , x0x1_subscript1_share2_wire , x0x2_subscript1_share2_wire , x0x3_subscript1_share2_wire , x0x4_subscript1_share2_wire , x0x5_subscript1_share2_wire , x0x6_subscript1_share2_wire , x0x7_subscript1_share2_wire , x1x2_subscript1_share2_wire , x1x3_subscript1_share2_wire , x1x4_subscript1_share2_wire , x1x5_subscript1_share2_wire , x1x6_subscript1_share2_wire , x1x7_subscript1_share2_wire , x2x3_subscript1_share2_wire , x2x4_subscript1_share2_wire , x2x5_subscript1_share2_wire , x2x6_subscript1_share2_wire , x2x7_subscript1_share2_wire , x3x4_subscript1_share2_wire , x3x5_subscript1_share2_wire , x3x6_subscript1_share2_wire , x3x7_subscript1_share2_wire , x4x5_subscript1_share2_wire , x4x6_subscript1_share2_wire , x4x7_subscript1_share2_wire , x5x6_subscript1_share2_wire , x5x7_subscript1_share2_wire , x6x7_subscript1_share2_wire , x0x1x2_subscript1_share2_wire , x0x1x3_subscript1_share2_wire , x0x1x4_subscript1_share2_wire , x0x1x5_subscript1_share2_wire , x0x1x6_subscript1_share2_wire , x0x1x7_subscript1_share2_wire , x0x2x3_subscript1_share2_wire , x0x2x4_subscript1_share2_wire , x0x2x5_subscript1_share2_wire , x0x2x6_subscript1_share2_wire , x0x2x7_subscript1_share2_wire , x0x3x4_subscript1_share2_wire , x0x3x5_subscript1_share2_wire , x0x3x6_subscript1_share2_wire , x0x3x7_subscript1_share2_wire , x0x4x5_subscript1_share2_wire , x0x4x6_subscript1_share2_wire , x0x4x7_subscript1_share2_wire , x0x5x6_subscript1_share2_wire , x0x5x7_subscript1_share2_wire , x0x6x7_subscript1_share2_wire , x1x2x3_subscript1_share2_wire , x1x2x4_subscript1_share2_wire , x1x2x5_subscript1_share2_wire , x1x2x6_subscript1_share2_wire , x1x2x7_subscript1_share2_wire , x1x3x4_subscript1_share2_wire , x1x3x5_subscript1_share2_wire , x1x3x6_subscript1_share2_wire , x1x3x7_subscript1_share2_wire , x1x4x5_subscript1_share2_wire , x1x4x6_subscript1_share2_wire , x1x4x7_subscript1_share2_wire , x1x5x6_subscript1_share2_wire , x1x5x7_subscript1_share2_wire , x1x6x7_subscript1_share2_wire , x2x3x4_subscript1_share2_wire , x2x3x5_subscript1_share2_wire , x2x3x6_subscript1_share2_wire , x2x3x7_subscript1_share2_wire , x2x4x5_subscript1_share2_wire , x2x4x6_subscript1_share2_wire , x2x4x7_subscript1_share2_wire , x2x5x6_subscript1_share2_wire , x2x5x7_subscript1_share2_wire , x2x6x7_subscript1_share2_wire , x3x4x5_subscript1_share2_wire , x3x4x6_subscript1_share2_wire , x3x4x7_subscript1_share2_wire , x3x5x6_subscript1_share2_wire , x3x5x7_subscript1_share2_wire , x3x6x7_subscript1_share2_wire , x4x5x6_subscript1_share2_wire , x4x5x7_subscript1_share2_wire , x4x6x7_subscript1_share2_wire , x5x6x7_subscript1_share2_wire , x0x1x2x3_subscript1_share2_wire , x0x1x2x4_subscript1_share2_wire , x0x1x2x5_subscript1_share2_wire , x0x1x2x6_subscript1_share2_wire , x0x1x2x7_subscript1_share2_wire , x0x1x3x4_subscript1_share2_wire , x0x1x3x5_subscript1_share2_wire , x0x1x3x6_subscript1_share2_wire , x0x1x3x7_subscript1_share2_wire , x0x1x4x5_subscript1_share2_wire , x0x1x4x6_subscript1_share2_wire , x0x1x4x7_subscript1_share2_wire , x0x1x5x6_subscript1_share2_wire , x0x1x5x7_subscript1_share2_wire , x0x1x6x7_subscript1_share2_wire , x0x2x3x4_subscript1_share2_wire , x0x2x3x5_subscript1_share2_wire , x0x2x3x6_subscript1_share2_wire , x0x2x3x7_subscript1_share2_wire , x0x2x4x5_subscript1_share2_wire , x0x2x4x6_subscript1_share2_wire , x0x2x4x7_subscript1_share2_wire , x0x2x5x6_subscript1_share2_wire , x0x2x5x7_subscript1_share2_wire , x0x2x6x7_subscript1_share2_wire , x0x3x4x5_subscript1_share2_wire , x0x3x4x6_subscript1_share2_wire , x0x3x4x7_subscript1_share2_wire , x0x3x5x6_subscript1_share2_wire , x0x3x5x7_subscript1_share2_wire , x0x3x6x7_subscript1_share2_wire , x0x4x5x6_subscript1_share2_wire , x0x4x5x7_subscript1_share2_wire , x0x4x6x7_subscript1_share2_wire , x0x5x6x7_subscript1_share2_wire , x1x2x3x4_subscript1_share2_wire , x1x2x3x5_subscript1_share2_wire , x1x2x3x6_subscript1_share2_wire , x1x2x3x7_subscript1_share2_wire , x1x2x4x5_subscript1_share2_wire , x1x2x4x6_subscript1_share2_wire , x1x2x4x7_subscript1_share2_wire , x1x2x5x6_subscript1_share2_wire , x1x2x5x7_subscript1_share2_wire , x1x2x6x7_subscript1_share2_wire , x1x3x4x5_subscript1_share2_wire , x1x3x4x6_subscript1_share2_wire , x1x3x4x7_subscript1_share2_wire , x1x3x5x6_subscript1_share2_wire , x1x3x5x7_subscript1_share2_wire , x1x3x6x7_subscript1_share2_wire , x1x4x5x6_subscript1_share2_wire , x1x4x5x7_subscript1_share2_wire , x1x4x6x7_subscript1_share2_wire , x1x5x6x7_subscript1_share2_wire , x2x3x4x5_subscript1_share2_wire , x2x3x4x6_subscript1_share2_wire , x2x3x4x7_subscript1_share2_wire , x2x3x5x6_subscript1_share2_wire , x2x3x5x7_subscript1_share2_wire , x2x3x6x7_subscript1_share2_wire , x2x4x5x6_subscript1_share2_wire , x2x4x5x7_subscript1_share2_wire , x2x4x6x7_subscript1_share2_wire , x2x5x6x7_subscript1_share2_wire , x3x4x5x6_subscript1_share2_wire , x3x4x5x7_subscript1_share2_wire , x3x4x6x7_subscript1_share2_wire , x3x5x6x7_subscript1_share2_wire , x4x5x6x7_subscript1_share2_wire , x0x1x2x3x4_subscript1_share2_wire , x0x1x2x3x5_subscript1_share2_wire , x0x1x2x3x6_subscript1_share2_wire , x0x1x2x3x7_subscript1_share2_wire , x0x1x2x4x5_subscript1_share2_wire , x0x1x2x4x6_subscript1_share2_wire , x0x1x2x4x7_subscript1_share2_wire , x0x1x2x5x6_subscript1_share2_wire , x0x1x2x5x7_subscript1_share2_wire , x0x1x2x6x7_subscript1_share2_wire , x0x1x3x4x5_subscript1_share2_wire , x0x1x3x4x6_subscript1_share2_wire , x0x1x3x4x7_subscript1_share2_wire , x0x1x3x5x6_subscript1_share2_wire , x0x1x3x5x7_subscript1_share2_wire , x0x1x3x6x7_subscript1_share2_wire , x0x1x4x5x6_subscript1_share2_wire , x0x1x4x5x7_subscript1_share2_wire , x0x1x4x6x7_subscript1_share2_wire , x0x1x5x6x7_subscript1_share2_wire , x0x2x3x4x5_subscript1_share2_wire , x0x2x3x4x6_subscript1_share2_wire , x0x2x3x4x7_subscript1_share2_wire , x0x2x3x5x6_subscript1_share2_wire , x0x2x3x5x7_subscript1_share2_wire , x0x2x3x6x7_subscript1_share2_wire , x0x2x4x5x6_subscript1_share2_wire , x0x2x4x5x7_subscript1_share2_wire , x0x2x4x6x7_subscript1_share2_wire , x0x2x5x6x7_subscript1_share2_wire , x0x3x4x5x6_subscript1_share2_wire , x0x3x4x5x7_subscript1_share2_wire , x0x3x4x6x7_subscript1_share2_wire , x0x3x5x6x7_subscript1_share2_wire , x0x4x5x6x7_subscript1_share2_wire , x1x2x3x4x5_subscript1_share2_wire , x1x2x3x4x6_subscript1_share2_wire , x1x2x3x4x7_subscript1_share2_wire , x1x2x3x5x6_subscript1_share2_wire , x1x2x3x5x7_subscript1_share2_wire , x1x2x3x6x7_subscript1_share2_wire , x1x2x4x5x6_subscript1_share2_wire , x1x2x4x5x7_subscript1_share2_wire , x1x2x4x6x7_subscript1_share2_wire , x1x2x5x6x7_subscript1_share2_wire , x1x3x4x5x6_subscript1_share2_wire , x1x3x4x5x7_subscript1_share2_wire , x1x3x4x6x7_subscript1_share2_wire , x1x3x5x6x7_subscript1_share2_wire , x1x4x5x6x7_subscript1_share2_wire , x2x3x4x5x6_subscript1_share2_wire , x2x3x4x5x7_subscript1_share2_wire , x2x3x4x6x7_subscript1_share2_wire , x2x3x5x6x7_subscript1_share2_wire , x2x4x5x6x7_subscript1_share2_wire , x3x4x5x6x7_subscript1_share2_wire , x0x1x2x3x4x5_subscript1_share2_wire , x0x1x2x3x4x6_subscript1_share2_wire , x0x1x2x3x4x7_subscript1_share2_wire , x0x1x2x3x5x6_subscript1_share2_wire , x0x1x2x3x5x7_subscript1_share2_wire , x0x1x2x3x6x7_subscript1_share2_wire , x0x1x2x4x5x6_subscript1_share2_wire , x0x1x2x4x5x7_subscript1_share2_wire , x0x1x2x4x6x7_subscript1_share2_wire , x0x1x2x5x6x7_subscript1_share2_wire , x0x1x3x4x5x6_subscript1_share2_wire , x0x1x3x4x5x7_subscript1_share2_wire , x0x1x3x4x6x7_subscript1_share2_wire , x0x1x3x5x6x7_subscript1_share2_wire , x0x1x4x5x6x7_subscript1_share2_wire , x0x2x3x4x5x6_subscript1_share2_wire , x0x2x3x4x5x7_subscript1_share2_wire , x0x2x3x4x6x7_subscript1_share2_wire , x0x2x3x5x6x7_subscript1_share2_wire , x0x2x4x5x6x7_subscript1_share2_wire , x0x3x4x5x6x7_subscript1_share2_wire , x1x2x3x4x5x6_subscript1_share2_wire , x1x2x3x4x5x7_subscript1_share2_wire , x1x2x3x4x6x7_subscript1_share2_wire , x1x2x3x5x6x7_subscript1_share2_wire , x1x2x4x5x6x7_subscript1_share2_wire , x1x3x4x5x6x7_subscript1_share2_wire , x2x3x4x5x6x7_subscript1_share2_wire , x0x1x2x3x4x5x6_subscript1_share2_wire , x0x1x2x3x4x5x7_subscript1_share2_wire , x0x1x2x3x4x6x7_subscript1_share2_wire , x0x1x2x3x5x6x7_subscript1_share2_wire , x0x1x2x4x5x6x7_subscript1_share2_wire , x0x1x3x4x5x6x7_subscript1_share2_wire , x0x2x3x4x5x6x7_subscript1_share2_wire , x1x2x3x4x5x6x7_subscript1_share2_wire ,
    x0_subscript1_share2_reg, x1_subscript1_share2_reg, x2_subscript1_share2_reg, x3_subscript1_share2_reg, x4_subscript1_share2_reg, x5_subscript1_share2_reg, x6_subscript1_share2_reg, x7_subscript1_share2_reg , x0x1_subscript1_share2_reg , x0x2_subscript1_share2_reg , x0x3_subscript1_share2_reg , x0x4_subscript1_share2_reg , x0x5_subscript1_share2_reg , x0x6_subscript1_share2_reg , x0x7_subscript1_share2_reg , x1x2_subscript1_share2_reg , x1x3_subscript1_share2_reg , x1x4_subscript1_share2_reg , x1x5_subscript1_share2_reg , x1x6_subscript1_share2_reg , x1x7_subscript1_share2_reg , x2x3_subscript1_share2_reg , x2x4_subscript1_share2_reg , x2x5_subscript1_share2_reg , x2x6_subscript1_share2_reg , x2x7_subscript1_share2_reg , x3x4_subscript1_share2_reg , x3x5_subscript1_share2_reg , x3x6_subscript1_share2_reg , x3x7_subscript1_share2_reg , x4x5_subscript1_share2_reg , x4x6_subscript1_share2_reg , x4x7_subscript1_share2_reg , x5x6_subscript1_share2_reg , x5x7_subscript1_share2_reg , x6x7_subscript1_share2_reg , x0x1x2_subscript1_share2_reg , x0x1x3_subscript1_share2_reg , x0x1x4_subscript1_share2_reg , x0x1x5_subscript1_share2_reg , x0x1x6_subscript1_share2_reg , x0x1x7_subscript1_share2_reg , x0x2x3_subscript1_share2_reg , x0x2x4_subscript1_share2_reg , x0x2x5_subscript1_share2_reg , x0x2x6_subscript1_share2_reg , x0x2x7_subscript1_share2_reg , x0x3x4_subscript1_share2_reg , x0x3x5_subscript1_share2_reg , x0x3x6_subscript1_share2_reg , x0x3x7_subscript1_share2_reg , x0x4x5_subscript1_share2_reg , x0x4x6_subscript1_share2_reg , x0x4x7_subscript1_share2_reg , x0x5x6_subscript1_share2_reg , x0x5x7_subscript1_share2_reg , x0x6x7_subscript1_share2_reg , x1x2x3_subscript1_share2_reg , x1x2x4_subscript1_share2_reg , x1x2x5_subscript1_share2_reg , x1x2x6_subscript1_share2_reg , x1x2x7_subscript1_share2_reg , x1x3x4_subscript1_share2_reg , x1x3x5_subscript1_share2_reg , x1x3x6_subscript1_share2_reg , x1x3x7_subscript1_share2_reg , x1x4x5_subscript1_share2_reg , x1x4x6_subscript1_share2_reg , x1x4x7_subscript1_share2_reg , x1x5x6_subscript1_share2_reg , x1x5x7_subscript1_share2_reg , x1x6x7_subscript1_share2_reg , x2x3x4_subscript1_share2_reg , x2x3x5_subscript1_share2_reg , x2x3x6_subscript1_share2_reg , x2x3x7_subscript1_share2_reg , x2x4x5_subscript1_share2_reg , x2x4x6_subscript1_share2_reg , x2x4x7_subscript1_share2_reg , x2x5x6_subscript1_share2_reg , x2x5x7_subscript1_share2_reg , x2x6x7_subscript1_share2_reg , x3x4x5_subscript1_share2_reg , x3x4x6_subscript1_share2_reg , x3x4x7_subscript1_share2_reg , x3x5x6_subscript1_share2_reg , x3x5x7_subscript1_share2_reg , x3x6x7_subscript1_share2_reg , x4x5x6_subscript1_share2_reg , x4x5x7_subscript1_share2_reg , x4x6x7_subscript1_share2_reg , x5x6x7_subscript1_share2_reg , x0x1x2x3_subscript1_share2_reg , x0x1x2x4_subscript1_share2_reg , x0x1x2x5_subscript1_share2_reg , x0x1x2x6_subscript1_share2_reg , x0x1x2x7_subscript1_share2_reg , x0x1x3x4_subscript1_share2_reg , x0x1x3x5_subscript1_share2_reg , x0x1x3x6_subscript1_share2_reg , x0x1x3x7_subscript1_share2_reg , x0x1x4x5_subscript1_share2_reg , x0x1x4x6_subscript1_share2_reg , x0x1x4x7_subscript1_share2_reg , x0x1x5x6_subscript1_share2_reg , x0x1x5x7_subscript1_share2_reg , x0x1x6x7_subscript1_share2_reg , x0x2x3x4_subscript1_share2_reg , x0x2x3x5_subscript1_share2_reg , x0x2x3x6_subscript1_share2_reg , x0x2x3x7_subscript1_share2_reg , x0x2x4x5_subscript1_share2_reg , x0x2x4x6_subscript1_share2_reg , x0x2x4x7_subscript1_share2_reg , x0x2x5x6_subscript1_share2_reg , x0x2x5x7_subscript1_share2_reg , x0x2x6x7_subscript1_share2_reg , x0x3x4x5_subscript1_share2_reg , x0x3x4x6_subscript1_share2_reg , x0x3x4x7_subscript1_share2_reg , x0x3x5x6_subscript1_share2_reg , x0x3x5x7_subscript1_share2_reg , x0x3x6x7_subscript1_share2_reg , x0x4x5x6_subscript1_share2_reg , x0x4x5x7_subscript1_share2_reg , x0x4x6x7_subscript1_share2_reg , x0x5x6x7_subscript1_share2_reg , x1x2x3x4_subscript1_share2_reg , x1x2x3x5_subscript1_share2_reg , x1x2x3x6_subscript1_share2_reg , x1x2x3x7_subscript1_share2_reg , x1x2x4x5_subscript1_share2_reg , x1x2x4x6_subscript1_share2_reg , x1x2x4x7_subscript1_share2_reg , x1x2x5x6_subscript1_share2_reg , x1x2x5x7_subscript1_share2_reg , x1x2x6x7_subscript1_share2_reg , x1x3x4x5_subscript1_share2_reg , x1x3x4x6_subscript1_share2_reg , x1x3x4x7_subscript1_share2_reg , x1x3x5x6_subscript1_share2_reg , x1x3x5x7_subscript1_share2_reg , x1x3x6x7_subscript1_share2_reg , x1x4x5x6_subscript1_share2_reg , x1x4x5x7_subscript1_share2_reg , x1x4x6x7_subscript1_share2_reg , x1x5x6x7_subscript1_share2_reg , x2x3x4x5_subscript1_share2_reg , x2x3x4x6_subscript1_share2_reg , x2x3x4x7_subscript1_share2_reg , x2x3x5x6_subscript1_share2_reg , x2x3x5x7_subscript1_share2_reg , x2x3x6x7_subscript1_share2_reg , x2x4x5x6_subscript1_share2_reg , x2x4x5x7_subscript1_share2_reg , x2x4x6x7_subscript1_share2_reg , x2x5x6x7_subscript1_share2_reg , x3x4x5x6_subscript1_share2_reg , x3x4x5x7_subscript1_share2_reg , x3x4x6x7_subscript1_share2_reg , x3x5x6x7_subscript1_share2_reg , x4x5x6x7_subscript1_share2_reg , x0x1x2x3x4_subscript1_share2_reg , x0x1x2x3x5_subscript1_share2_reg , x0x1x2x3x6_subscript1_share2_reg , x0x1x2x3x7_subscript1_share2_reg , x0x1x2x4x5_subscript1_share2_reg , x0x1x2x4x6_subscript1_share2_reg , x0x1x2x4x7_subscript1_share2_reg , x0x1x2x5x6_subscript1_share2_reg , x0x1x2x5x7_subscript1_share2_reg , x0x1x2x6x7_subscript1_share2_reg , x0x1x3x4x5_subscript1_share2_reg , x0x1x3x4x6_subscript1_share2_reg , x0x1x3x4x7_subscript1_share2_reg , x0x1x3x5x6_subscript1_share2_reg , x0x1x3x5x7_subscript1_share2_reg , x0x1x3x6x7_subscript1_share2_reg , x0x1x4x5x6_subscript1_share2_reg , x0x1x4x5x7_subscript1_share2_reg , x0x1x4x6x7_subscript1_share2_reg , x0x1x5x6x7_subscript1_share2_reg , x0x2x3x4x5_subscript1_share2_reg , x0x2x3x4x6_subscript1_share2_reg , x0x2x3x4x7_subscript1_share2_reg , x0x2x3x5x6_subscript1_share2_reg , x0x2x3x5x7_subscript1_share2_reg , x0x2x3x6x7_subscript1_share2_reg , x0x2x4x5x6_subscript1_share2_reg , x0x2x4x5x7_subscript1_share2_reg , x0x2x4x6x7_subscript1_share2_reg , x0x2x5x6x7_subscript1_share2_reg , x0x3x4x5x6_subscript1_share2_reg , x0x3x4x5x7_subscript1_share2_reg , x0x3x4x6x7_subscript1_share2_reg , x0x3x5x6x7_subscript1_share2_reg , x0x4x5x6x7_subscript1_share2_reg , x1x2x3x4x5_subscript1_share2_reg , x1x2x3x4x6_subscript1_share2_reg , x1x2x3x4x7_subscript1_share2_reg , x1x2x3x5x6_subscript1_share2_reg , x1x2x3x5x7_subscript1_share2_reg , x1x2x3x6x7_subscript1_share2_reg , x1x2x4x5x6_subscript1_share2_reg , x1x2x4x5x7_subscript1_share2_reg , x1x2x4x6x7_subscript1_share2_reg , x1x2x5x6x7_subscript1_share2_reg , x1x3x4x5x6_subscript1_share2_reg , x1x3x4x5x7_subscript1_share2_reg , x1x3x4x6x7_subscript1_share2_reg , x1x3x5x6x7_subscript1_share2_reg , x1x4x5x6x7_subscript1_share2_reg , x2x3x4x5x6_subscript1_share2_reg , x2x3x4x5x7_subscript1_share2_reg , x2x3x4x6x7_subscript1_share2_reg , x2x3x5x6x7_subscript1_share2_reg , x2x4x5x6x7_subscript1_share2_reg , x3x4x5x6x7_subscript1_share2_reg , x0x1x2x3x4x5_subscript1_share2_reg , x0x1x2x3x4x6_subscript1_share2_reg , x0x1x2x3x4x7_subscript1_share2_reg , x0x1x2x3x5x6_subscript1_share2_reg , x0x1x2x3x5x7_subscript1_share2_reg , x0x1x2x3x6x7_subscript1_share2_reg , x0x1x2x4x5x6_subscript1_share2_reg , x0x1x2x4x5x7_subscript1_share2_reg , x0x1x2x4x6x7_subscript1_share2_reg , x0x1x2x5x6x7_subscript1_share2_reg , x0x1x3x4x5x6_subscript1_share2_reg , x0x1x3x4x5x7_subscript1_share2_reg , x0x1x3x4x6x7_subscript1_share2_reg , x0x1x3x5x6x7_subscript1_share2_reg , x0x1x4x5x6x7_subscript1_share2_reg , x0x2x3x4x5x6_subscript1_share2_reg , x0x2x3x4x5x7_subscript1_share2_reg , x0x2x3x4x6x7_subscript1_share2_reg , x0x2x3x5x6x7_subscript1_share2_reg , x0x2x4x5x6x7_subscript1_share2_reg , x0x3x4x5x6x7_subscript1_share2_reg , x1x2x3x4x5x6_subscript1_share2_reg , x1x2x3x4x5x7_subscript1_share2_reg , x1x2x3x4x6x7_subscript1_share2_reg , x1x2x3x5x6x7_subscript1_share2_reg , x1x2x4x5x6x7_subscript1_share2_reg , x1x3x4x5x6x7_subscript1_share2_reg , x2x3x4x5x6x7_subscript1_share2_reg , x0x1x2x3x4x5x6_subscript1_share2_reg , x0x1x2x3x4x5x7_subscript1_share2_reg , x0x1x2x3x4x6x7_subscript1_share2_reg , x0x1x2x3x5x6x7_subscript1_share2_reg , x0x1x2x4x5x6x7_subscript1_share2_reg , x0x1x3x4x5x6x7_subscript1_share2_reg , x0x2x3x4x5x6x7_subscript1_share2_reg , x1x2x3x4x5x6x7_subscript1_share2_reg 
);
register_array_AES_oneshare second_cycle_share3_reg (
    clk,
    x0_subscript1_share3_wire, x1_subscript1_share3_wire, x2_subscript1_share3_wire, x3_subscript1_share3_wire, x4_subscript1_share3_wire, x5_subscript1_share3_wire, x6_subscript1_share3_wire, x7_subscript1_share3_wire , x0x1_subscript1_share3_wire , x0x2_subscript1_share3_wire , x0x3_subscript1_share3_wire , x0x4_subscript1_share3_wire , x0x5_subscript1_share3_wire , x0x6_subscript1_share3_wire , x0x7_subscript1_share3_wire , x1x2_subscript1_share3_wire , x1x3_subscript1_share3_wire , x1x4_subscript1_share3_wire , x1x5_subscript1_share3_wire , x1x6_subscript1_share3_wire , x1x7_subscript1_share3_wire , x2x3_subscript1_share3_wire , x2x4_subscript1_share3_wire , x2x5_subscript1_share3_wire , x2x6_subscript1_share3_wire , x2x7_subscript1_share3_wire , x3x4_subscript1_share3_wire , x3x5_subscript1_share3_wire , x3x6_subscript1_share3_wire , x3x7_subscript1_share3_wire , x4x5_subscript1_share3_wire , x4x6_subscript1_share3_wire , x4x7_subscript1_share3_wire , x5x6_subscript1_share3_wire , x5x7_subscript1_share3_wire , x6x7_subscript1_share3_wire , x0x1x2_subscript1_share3_wire , x0x1x3_subscript1_share3_wire , x0x1x4_subscript1_share3_wire , x0x1x5_subscript1_share3_wire , x0x1x6_subscript1_share3_wire , x0x1x7_subscript1_share3_wire , x0x2x3_subscript1_share3_wire , x0x2x4_subscript1_share3_wire , x0x2x5_subscript1_share3_wire , x0x2x6_subscript1_share3_wire , x0x2x7_subscript1_share3_wire , x0x3x4_subscript1_share3_wire , x0x3x5_subscript1_share3_wire , x0x3x6_subscript1_share3_wire , x0x3x7_subscript1_share3_wire , x0x4x5_subscript1_share3_wire , x0x4x6_subscript1_share3_wire , x0x4x7_subscript1_share3_wire , x0x5x6_subscript1_share3_wire , x0x5x7_subscript1_share3_wire , x0x6x7_subscript1_share3_wire , x1x2x3_subscript1_share3_wire , x1x2x4_subscript1_share3_wire , x1x2x5_subscript1_share3_wire , x1x2x6_subscript1_share3_wire , x1x2x7_subscript1_share3_wire , x1x3x4_subscript1_share3_wire , x1x3x5_subscript1_share3_wire , x1x3x6_subscript1_share3_wire , x1x3x7_subscript1_share3_wire , x1x4x5_subscript1_share3_wire , x1x4x6_subscript1_share3_wire , x1x4x7_subscript1_share3_wire , x1x5x6_subscript1_share3_wire , x1x5x7_subscript1_share3_wire , x1x6x7_subscript1_share3_wire , x2x3x4_subscript1_share3_wire , x2x3x5_subscript1_share3_wire , x2x3x6_subscript1_share3_wire , x2x3x7_subscript1_share3_wire , x2x4x5_subscript1_share3_wire , x2x4x6_subscript1_share3_wire , x2x4x7_subscript1_share3_wire , x2x5x6_subscript1_share3_wire , x2x5x7_subscript1_share3_wire , x2x6x7_subscript1_share3_wire , x3x4x5_subscript1_share3_wire , x3x4x6_subscript1_share3_wire , x3x4x7_subscript1_share3_wire , x3x5x6_subscript1_share3_wire , x3x5x7_subscript1_share3_wire , x3x6x7_subscript1_share3_wire , x4x5x6_subscript1_share3_wire , x4x5x7_subscript1_share3_wire , x4x6x7_subscript1_share3_wire , x5x6x7_subscript1_share3_wire , x0x1x2x3_subscript1_share3_wire , x0x1x2x4_subscript1_share3_wire , x0x1x2x5_subscript1_share3_wire , x0x1x2x6_subscript1_share3_wire , x0x1x2x7_subscript1_share3_wire , x0x1x3x4_subscript1_share3_wire , x0x1x3x5_subscript1_share3_wire , x0x1x3x6_subscript1_share3_wire , x0x1x3x7_subscript1_share3_wire , x0x1x4x5_subscript1_share3_wire , x0x1x4x6_subscript1_share3_wire , x0x1x4x7_subscript1_share3_wire , x0x1x5x6_subscript1_share3_wire , x0x1x5x7_subscript1_share3_wire , x0x1x6x7_subscript1_share3_wire , x0x2x3x4_subscript1_share3_wire , x0x2x3x5_subscript1_share3_wire , x0x2x3x6_subscript1_share3_wire , x0x2x3x7_subscript1_share3_wire , x0x2x4x5_subscript1_share3_wire , x0x2x4x6_subscript1_share3_wire , x0x2x4x7_subscript1_share3_wire , x0x2x5x6_subscript1_share3_wire , x0x2x5x7_subscript1_share3_wire , x0x2x6x7_subscript1_share3_wire , x0x3x4x5_subscript1_share3_wire , x0x3x4x6_subscript1_share3_wire , x0x3x4x7_subscript1_share3_wire , x0x3x5x6_subscript1_share3_wire , x0x3x5x7_subscript1_share3_wire , x0x3x6x7_subscript1_share3_wire , x0x4x5x6_subscript1_share3_wire , x0x4x5x7_subscript1_share3_wire , x0x4x6x7_subscript1_share3_wire , x0x5x6x7_subscript1_share3_wire , x1x2x3x4_subscript1_share3_wire , x1x2x3x5_subscript1_share3_wire , x1x2x3x6_subscript1_share3_wire , x1x2x3x7_subscript1_share3_wire , x1x2x4x5_subscript1_share3_wire , x1x2x4x6_subscript1_share3_wire , x1x2x4x7_subscript1_share3_wire , x1x2x5x6_subscript1_share3_wire , x1x2x5x7_subscript1_share3_wire , x1x2x6x7_subscript1_share3_wire , x1x3x4x5_subscript1_share3_wire , x1x3x4x6_subscript1_share3_wire , x1x3x4x7_subscript1_share3_wire , x1x3x5x6_subscript1_share3_wire , x1x3x5x7_subscript1_share3_wire , x1x3x6x7_subscript1_share3_wire , x1x4x5x6_subscript1_share3_wire , x1x4x5x7_subscript1_share3_wire , x1x4x6x7_subscript1_share3_wire , x1x5x6x7_subscript1_share3_wire , x2x3x4x5_subscript1_share3_wire , x2x3x4x6_subscript1_share3_wire , x2x3x4x7_subscript1_share3_wire , x2x3x5x6_subscript1_share3_wire , x2x3x5x7_subscript1_share3_wire , x2x3x6x7_subscript1_share3_wire , x2x4x5x6_subscript1_share3_wire , x2x4x5x7_subscript1_share3_wire , x2x4x6x7_subscript1_share3_wire , x2x5x6x7_subscript1_share3_wire , x3x4x5x6_subscript1_share3_wire , x3x4x5x7_subscript1_share3_wire , x3x4x6x7_subscript1_share3_wire , x3x5x6x7_subscript1_share3_wire , x4x5x6x7_subscript1_share3_wire , x0x1x2x3x4_subscript1_share3_wire , x0x1x2x3x5_subscript1_share3_wire , x0x1x2x3x6_subscript1_share3_wire , x0x1x2x3x7_subscript1_share3_wire , x0x1x2x4x5_subscript1_share3_wire , x0x1x2x4x6_subscript1_share3_wire , x0x1x2x4x7_subscript1_share3_wire , x0x1x2x5x6_subscript1_share3_wire , x0x1x2x5x7_subscript1_share3_wire , x0x1x2x6x7_subscript1_share3_wire , x0x1x3x4x5_subscript1_share3_wire , x0x1x3x4x6_subscript1_share3_wire , x0x1x3x4x7_subscript1_share3_wire , x0x1x3x5x6_subscript1_share3_wire , x0x1x3x5x7_subscript1_share3_wire , x0x1x3x6x7_subscript1_share3_wire , x0x1x4x5x6_subscript1_share3_wire , x0x1x4x5x7_subscript1_share3_wire , x0x1x4x6x7_subscript1_share3_wire , x0x1x5x6x7_subscript1_share3_wire , x0x2x3x4x5_subscript1_share3_wire , x0x2x3x4x6_subscript1_share3_wire , x0x2x3x4x7_subscript1_share3_wire , x0x2x3x5x6_subscript1_share3_wire , x0x2x3x5x7_subscript1_share3_wire , x0x2x3x6x7_subscript1_share3_wire , x0x2x4x5x6_subscript1_share3_wire , x0x2x4x5x7_subscript1_share3_wire , x0x2x4x6x7_subscript1_share3_wire , x0x2x5x6x7_subscript1_share3_wire , x0x3x4x5x6_subscript1_share3_wire , x0x3x4x5x7_subscript1_share3_wire , x0x3x4x6x7_subscript1_share3_wire , x0x3x5x6x7_subscript1_share3_wire , x0x4x5x6x7_subscript1_share3_wire , x1x2x3x4x5_subscript1_share3_wire , x1x2x3x4x6_subscript1_share3_wire , x1x2x3x4x7_subscript1_share3_wire , x1x2x3x5x6_subscript1_share3_wire , x1x2x3x5x7_subscript1_share3_wire , x1x2x3x6x7_subscript1_share3_wire , x1x2x4x5x6_subscript1_share3_wire , x1x2x4x5x7_subscript1_share3_wire , x1x2x4x6x7_subscript1_share3_wire , x1x2x5x6x7_subscript1_share3_wire , x1x3x4x5x6_subscript1_share3_wire , x1x3x4x5x7_subscript1_share3_wire , x1x3x4x6x7_subscript1_share3_wire , x1x3x5x6x7_subscript1_share3_wire , x1x4x5x6x7_subscript1_share3_wire , x2x3x4x5x6_subscript1_share3_wire , x2x3x4x5x7_subscript1_share3_wire , x2x3x4x6x7_subscript1_share3_wire , x2x3x5x6x7_subscript1_share3_wire , x2x4x5x6x7_subscript1_share3_wire , x3x4x5x6x7_subscript1_share3_wire , x0x1x2x3x4x5_subscript1_share3_wire , x0x1x2x3x4x6_subscript1_share3_wire , x0x1x2x3x4x7_subscript1_share3_wire , x0x1x2x3x5x6_subscript1_share3_wire , x0x1x2x3x5x7_subscript1_share3_wire , x0x1x2x3x6x7_subscript1_share3_wire , x0x1x2x4x5x6_subscript1_share3_wire , x0x1x2x4x5x7_subscript1_share3_wire , x0x1x2x4x6x7_subscript1_share3_wire , x0x1x2x5x6x7_subscript1_share3_wire , x0x1x3x4x5x6_subscript1_share3_wire , x0x1x3x4x5x7_subscript1_share3_wire , x0x1x3x4x6x7_subscript1_share3_wire , x0x1x3x5x6x7_subscript1_share3_wire , x0x1x4x5x6x7_subscript1_share3_wire , x0x2x3x4x5x6_subscript1_share3_wire , x0x2x3x4x5x7_subscript1_share3_wire , x0x2x3x4x6x7_subscript1_share3_wire , x0x2x3x5x6x7_subscript1_share3_wire , x0x2x4x5x6x7_subscript1_share3_wire , x0x3x4x5x6x7_subscript1_share3_wire , x1x2x3x4x5x6_subscript1_share3_wire , x1x2x3x4x5x7_subscript1_share3_wire , x1x2x3x4x6x7_subscript1_share3_wire , x1x2x3x5x6x7_subscript1_share3_wire , x1x2x4x5x6x7_subscript1_share3_wire , x1x3x4x5x6x7_subscript1_share3_wire , x2x3x4x5x6x7_subscript1_share3_wire , x0x1x2x3x4x5x6_subscript1_share3_wire , x0x1x2x3x4x5x7_subscript1_share3_wire , x0x1x2x3x4x6x7_subscript1_share3_wire , x0x1x2x3x5x6x7_subscript1_share3_wire , x0x1x2x4x5x6x7_subscript1_share3_wire , x0x1x3x4x5x6x7_subscript1_share3_wire , x0x2x3x4x5x6x7_subscript1_share3_wire , x1x2x3x4x5x6x7_subscript1_share3_wire ,
    x0_subscript1_share3_reg, x1_subscript1_share3_reg, x2_subscript1_share3_reg, x3_subscript1_share3_reg, x4_subscript1_share3_reg, x5_subscript1_share3_reg, x6_subscript1_share3_reg, x7_subscript1_share3_reg , x0x1_subscript1_share3_reg , x0x2_subscript1_share3_reg , x0x3_subscript1_share3_reg , x0x4_subscript1_share3_reg , x0x5_subscript1_share3_reg , x0x6_subscript1_share3_reg , x0x7_subscript1_share3_reg , x1x2_subscript1_share3_reg , x1x3_subscript1_share3_reg , x1x4_subscript1_share3_reg , x1x5_subscript1_share3_reg , x1x6_subscript1_share3_reg , x1x7_subscript1_share3_reg , x2x3_subscript1_share3_reg , x2x4_subscript1_share3_reg , x2x5_subscript1_share3_reg , x2x6_subscript1_share3_reg , x2x7_subscript1_share3_reg , x3x4_subscript1_share3_reg , x3x5_subscript1_share3_reg , x3x6_subscript1_share3_reg , x3x7_subscript1_share3_reg , x4x5_subscript1_share3_reg , x4x6_subscript1_share3_reg , x4x7_subscript1_share3_reg , x5x6_subscript1_share3_reg , x5x7_subscript1_share3_reg , x6x7_subscript1_share3_reg , x0x1x2_subscript1_share3_reg , x0x1x3_subscript1_share3_reg , x0x1x4_subscript1_share3_reg , x0x1x5_subscript1_share3_reg , x0x1x6_subscript1_share3_reg , x0x1x7_subscript1_share3_reg , x0x2x3_subscript1_share3_reg , x0x2x4_subscript1_share3_reg , x0x2x5_subscript1_share3_reg , x0x2x6_subscript1_share3_reg , x0x2x7_subscript1_share3_reg , x0x3x4_subscript1_share3_reg , x0x3x5_subscript1_share3_reg , x0x3x6_subscript1_share3_reg , x0x3x7_subscript1_share3_reg , x0x4x5_subscript1_share3_reg , x0x4x6_subscript1_share3_reg , x0x4x7_subscript1_share3_reg , x0x5x6_subscript1_share3_reg , x0x5x7_subscript1_share3_reg , x0x6x7_subscript1_share3_reg , x1x2x3_subscript1_share3_reg , x1x2x4_subscript1_share3_reg , x1x2x5_subscript1_share3_reg , x1x2x6_subscript1_share3_reg , x1x2x7_subscript1_share3_reg , x1x3x4_subscript1_share3_reg , x1x3x5_subscript1_share3_reg , x1x3x6_subscript1_share3_reg , x1x3x7_subscript1_share3_reg , x1x4x5_subscript1_share3_reg , x1x4x6_subscript1_share3_reg , x1x4x7_subscript1_share3_reg , x1x5x6_subscript1_share3_reg , x1x5x7_subscript1_share3_reg , x1x6x7_subscript1_share3_reg , x2x3x4_subscript1_share3_reg , x2x3x5_subscript1_share3_reg , x2x3x6_subscript1_share3_reg , x2x3x7_subscript1_share3_reg , x2x4x5_subscript1_share3_reg , x2x4x6_subscript1_share3_reg , x2x4x7_subscript1_share3_reg , x2x5x6_subscript1_share3_reg , x2x5x7_subscript1_share3_reg , x2x6x7_subscript1_share3_reg , x3x4x5_subscript1_share3_reg , x3x4x6_subscript1_share3_reg , x3x4x7_subscript1_share3_reg , x3x5x6_subscript1_share3_reg , x3x5x7_subscript1_share3_reg , x3x6x7_subscript1_share3_reg , x4x5x6_subscript1_share3_reg , x4x5x7_subscript1_share3_reg , x4x6x7_subscript1_share3_reg , x5x6x7_subscript1_share3_reg , x0x1x2x3_subscript1_share3_reg , x0x1x2x4_subscript1_share3_reg , x0x1x2x5_subscript1_share3_reg , x0x1x2x6_subscript1_share3_reg , x0x1x2x7_subscript1_share3_reg , x0x1x3x4_subscript1_share3_reg , x0x1x3x5_subscript1_share3_reg , x0x1x3x6_subscript1_share3_reg , x0x1x3x7_subscript1_share3_reg , x0x1x4x5_subscript1_share3_reg , x0x1x4x6_subscript1_share3_reg , x0x1x4x7_subscript1_share3_reg , x0x1x5x6_subscript1_share3_reg , x0x1x5x7_subscript1_share3_reg , x0x1x6x7_subscript1_share3_reg , x0x2x3x4_subscript1_share3_reg , x0x2x3x5_subscript1_share3_reg , x0x2x3x6_subscript1_share3_reg , x0x2x3x7_subscript1_share3_reg , x0x2x4x5_subscript1_share3_reg , x0x2x4x6_subscript1_share3_reg , x0x2x4x7_subscript1_share3_reg , x0x2x5x6_subscript1_share3_reg , x0x2x5x7_subscript1_share3_reg , x0x2x6x7_subscript1_share3_reg , x0x3x4x5_subscript1_share3_reg , x0x3x4x6_subscript1_share3_reg , x0x3x4x7_subscript1_share3_reg , x0x3x5x6_subscript1_share3_reg , x0x3x5x7_subscript1_share3_reg , x0x3x6x7_subscript1_share3_reg , x0x4x5x6_subscript1_share3_reg , x0x4x5x7_subscript1_share3_reg , x0x4x6x7_subscript1_share3_reg , x0x5x6x7_subscript1_share3_reg , x1x2x3x4_subscript1_share3_reg , x1x2x3x5_subscript1_share3_reg , x1x2x3x6_subscript1_share3_reg , x1x2x3x7_subscript1_share3_reg , x1x2x4x5_subscript1_share3_reg , x1x2x4x6_subscript1_share3_reg , x1x2x4x7_subscript1_share3_reg , x1x2x5x6_subscript1_share3_reg , x1x2x5x7_subscript1_share3_reg , x1x2x6x7_subscript1_share3_reg , x1x3x4x5_subscript1_share3_reg , x1x3x4x6_subscript1_share3_reg , x1x3x4x7_subscript1_share3_reg , x1x3x5x6_subscript1_share3_reg , x1x3x5x7_subscript1_share3_reg , x1x3x6x7_subscript1_share3_reg , x1x4x5x6_subscript1_share3_reg , x1x4x5x7_subscript1_share3_reg , x1x4x6x7_subscript1_share3_reg , x1x5x6x7_subscript1_share3_reg , x2x3x4x5_subscript1_share3_reg , x2x3x4x6_subscript1_share3_reg , x2x3x4x7_subscript1_share3_reg , x2x3x5x6_subscript1_share3_reg , x2x3x5x7_subscript1_share3_reg , x2x3x6x7_subscript1_share3_reg , x2x4x5x6_subscript1_share3_reg , x2x4x5x7_subscript1_share3_reg , x2x4x6x7_subscript1_share3_reg , x2x5x6x7_subscript1_share3_reg , x3x4x5x6_subscript1_share3_reg , x3x4x5x7_subscript1_share3_reg , x3x4x6x7_subscript1_share3_reg , x3x5x6x7_subscript1_share3_reg , x4x5x6x7_subscript1_share3_reg , x0x1x2x3x4_subscript1_share3_reg , x0x1x2x3x5_subscript1_share3_reg , x0x1x2x3x6_subscript1_share3_reg , x0x1x2x3x7_subscript1_share3_reg , x0x1x2x4x5_subscript1_share3_reg , x0x1x2x4x6_subscript1_share3_reg , x0x1x2x4x7_subscript1_share3_reg , x0x1x2x5x6_subscript1_share3_reg , x0x1x2x5x7_subscript1_share3_reg , x0x1x2x6x7_subscript1_share3_reg , x0x1x3x4x5_subscript1_share3_reg , x0x1x3x4x6_subscript1_share3_reg , x0x1x3x4x7_subscript1_share3_reg , x0x1x3x5x6_subscript1_share3_reg , x0x1x3x5x7_subscript1_share3_reg , x0x1x3x6x7_subscript1_share3_reg , x0x1x4x5x6_subscript1_share3_reg , x0x1x4x5x7_subscript1_share3_reg , x0x1x4x6x7_subscript1_share3_reg , x0x1x5x6x7_subscript1_share3_reg , x0x2x3x4x5_subscript1_share3_reg , x0x2x3x4x6_subscript1_share3_reg , x0x2x3x4x7_subscript1_share3_reg , x0x2x3x5x6_subscript1_share3_reg , x0x2x3x5x7_subscript1_share3_reg , x0x2x3x6x7_subscript1_share3_reg , x0x2x4x5x6_subscript1_share3_reg , x0x2x4x5x7_subscript1_share3_reg , x0x2x4x6x7_subscript1_share3_reg , x0x2x5x6x7_subscript1_share3_reg , x0x3x4x5x6_subscript1_share3_reg , x0x3x4x5x7_subscript1_share3_reg , x0x3x4x6x7_subscript1_share3_reg , x0x3x5x6x7_subscript1_share3_reg , x0x4x5x6x7_subscript1_share3_reg , x1x2x3x4x5_subscript1_share3_reg , x1x2x3x4x6_subscript1_share3_reg , x1x2x3x4x7_subscript1_share3_reg , x1x2x3x5x6_subscript1_share3_reg , x1x2x3x5x7_subscript1_share3_reg , x1x2x3x6x7_subscript1_share3_reg , x1x2x4x5x6_subscript1_share3_reg , x1x2x4x5x7_subscript1_share3_reg , x1x2x4x6x7_subscript1_share3_reg , x1x2x5x6x7_subscript1_share3_reg , x1x3x4x5x6_subscript1_share3_reg , x1x3x4x5x7_subscript1_share3_reg , x1x3x4x6x7_subscript1_share3_reg , x1x3x5x6x7_subscript1_share3_reg , x1x4x5x6x7_subscript1_share3_reg , x2x3x4x5x6_subscript1_share3_reg , x2x3x4x5x7_subscript1_share3_reg , x2x3x4x6x7_subscript1_share3_reg , x2x3x5x6x7_subscript1_share3_reg , x2x4x5x6x7_subscript1_share3_reg , x3x4x5x6x7_subscript1_share3_reg , x0x1x2x3x4x5_subscript1_share3_reg , x0x1x2x3x4x6_subscript1_share3_reg , x0x1x2x3x4x7_subscript1_share3_reg , x0x1x2x3x5x6_subscript1_share3_reg , x0x1x2x3x5x7_subscript1_share3_reg , x0x1x2x3x6x7_subscript1_share3_reg , x0x1x2x4x5x6_subscript1_share3_reg , x0x1x2x4x5x7_subscript1_share3_reg , x0x1x2x4x6x7_subscript1_share3_reg , x0x1x2x5x6x7_subscript1_share3_reg , x0x1x3x4x5x6_subscript1_share3_reg , x0x1x3x4x5x7_subscript1_share3_reg , x0x1x3x4x6x7_subscript1_share3_reg , x0x1x3x5x6x7_subscript1_share3_reg , x0x1x4x5x6x7_subscript1_share3_reg , x0x2x3x4x5x6_subscript1_share3_reg , x0x2x3x4x5x7_subscript1_share3_reg , x0x2x3x4x6x7_subscript1_share3_reg , x0x2x3x5x6x7_subscript1_share3_reg , x0x2x4x5x6x7_subscript1_share3_reg , x0x3x4x5x6x7_subscript1_share3_reg , x1x2x3x4x5x6_subscript1_share3_reg , x1x2x3x4x5x7_subscript1_share3_reg , x1x2x3x4x6x7_subscript1_share3_reg , x1x2x3x5x6x7_subscript1_share3_reg , x1x2x4x5x6x7_subscript1_share3_reg , x1x3x4x5x6x7_subscript1_share3_reg , x2x3x4x5x6x7_subscript1_share3_reg , x0x1x2x3x4x5x6_subscript1_share3_reg , x0x1x2x3x4x5x7_subscript1_share3_reg , x0x1x2x3x4x6x7_subscript1_share3_reg , x0x1x2x3x5x6x7_subscript1_share3_reg , x0x1x2x4x5x6x7_subscript1_share3_reg , x0x1x3x4x5x6x7_subscript1_share3_reg , x0x2x3x4x5x6x7_subscript1_share3_reg , x1x2x3x4x5x6x7_subscript1_share3_reg 
);

register_array_8bit_AES  reg_second_cycle_pipeline_share3 (clk , x0_pipelined_share3_reg, x1_pipelined_share3_reg, x2_pipelined_share3_reg, x3_pipelined_share3_reg, x4_pipelined_share3_reg, x5_pipelined_share3_reg, x6_pipelined_share3_reg, x7_pipelined_share3_reg, x0_pipelined2_share3_reg, x1_pipelined2_share3_reg, x2_pipelined2_share3_reg, x3_pipelined2_share3_reg, x4_pipelined2_share3_reg, x5_pipelined2_share3_reg, x6_pipelined2_share3_reg, x7_pipelined2_share3_reg );



// Cycle 3

wire sbox_out1_share1, sbox_out2_share1, sbox_out3_share1, sbox_out4_share1, sbox_out5_share1, sbox_out6_share1, sbox_out7_share1, sbox_out8_share1 ;
wire sbox_out1_share2, sbox_out2_share2, sbox_out3_share2, sbox_out4_share2, sbox_out5_share2, sbox_out6_share2, sbox_out7_share2, sbox_out8_share2 ;
wire sbox_out1_share3, sbox_out2_share3, sbox_out3_share3, sbox_out4_share3, sbox_out5_share3, sbox_out6_share3, sbox_out7_share3, sbox_out8_share3 ;


combi_logic_cycle3_output_share1 inst_cycle3_share1 (
    x0_subscript1_share1_reg , x2_subscript1_share1_reg , x3_subscript1_share1_reg , x4_subscript1_share1_reg , x6_subscript1_share1_reg , x7_subscript1_share1_reg , x1_subscript1_share1_reg , x5_subscript1_share1_reg , x0x1_subscript1_share1_reg , x0x4_subscript1_share1_reg , x0x5_subscript1_share1_reg , x0x6_subscript1_share1_reg , x1x2_subscript1_share1_reg , x1x3_subscript1_share1_reg , x1x4_subscript1_share1_reg , x1x6_subscript1_share1_reg , x2x3_subscript1_share1_reg , x2x4_subscript1_share1_reg , x2x6_subscript1_share1_reg , x2x7_subscript1_share1_reg , x4x6_subscript1_share1_reg , x5x6_subscript1_share1_reg , x5x7_subscript1_share1_reg , x6x7_subscript1_share1_reg , x0x2_subscript1_share1_reg , x0x3_subscript1_share1_reg , x0x7_subscript1_share1_reg , x1x7_subscript1_share1_reg , x3x7_subscript1_share1_reg , x4x5_subscript1_share1_reg , x3x4_subscript1_share1_reg , x4x7_subscript1_share1_reg , x3x6_subscript1_share1_reg , x1x5_subscript1_share1_reg , x2x5_subscript1_share1_reg , x3x5_subscript1_share1_reg , x0x1x4_subscript1_share1_reg , x0x1x6_subscript1_share1_reg , x0x1x7_subscript1_share1_reg , x0x2x4_subscript1_share1_reg , x0x2x5_subscript1_share1_reg , x0x2x6_subscript1_share1_reg , x0x2x7_subscript1_share1_reg , x0x3x4_subscript1_share1_reg , x0x3x5_subscript1_share1_reg , x0x3x6_subscript1_share1_reg , x0x4x6_subscript1_share1_reg , x0x4x7_subscript1_share1_reg , x1x2x3_subscript1_share1_reg , x1x2x4_subscript1_share1_reg , x1x2x6_subscript1_share1_reg , x1x3x4_subscript1_share1_reg , x1x3x7_subscript1_share1_reg , x1x4x6_subscript1_share1_reg , x1x5x6_subscript1_share1_reg , x2x3x5_subscript1_share1_reg , x2x3x7_subscript1_share1_reg , x2x4x7_subscript1_share1_reg , x2x5x6_subscript1_share1_reg , x2x5x7_subscript1_share1_reg , x2x6x7_subscript1_share1_reg , x3x4x7_subscript1_share1_reg , x3x5x7_subscript1_share1_reg , x3x6x7_subscript1_share1_reg , x4x5x6_subscript1_share1_reg , x5x6x7_subscript1_share1_reg , x0x1x3_subscript1_share1_reg , x0x2x3_subscript1_share1_reg , x0x4x5_subscript1_share1_reg , x0x5x7_subscript1_share1_reg , x0x6x7_subscript1_share1_reg , x1x3x5_subscript1_share1_reg , x1x3x6_subscript1_share1_reg , x1x4x7_subscript1_share1_reg , x2x3x4_subscript1_share1_reg , x2x3x6_subscript1_share1_reg , x3x4x6_subscript1_share1_reg , x3x5x6_subscript1_share1_reg , x0x1x5_subscript1_share1_reg , x0x3x7_subscript1_share1_reg , x1x2x5_subscript1_share1_reg , x1x2x7_subscript1_share1_reg , x1x4x5_subscript1_share1_reg , x1x5x7_subscript1_share1_reg , x2x4x5_subscript1_share1_reg , x3x4x5_subscript1_share1_reg , x4x6x7_subscript1_share1_reg , x1x6x7_subscript1_share1_reg , x4x5x7_subscript1_share1_reg , x0x1x2_subscript1_share1_reg , x0x5x6_subscript1_share1_reg , x2x4x6_subscript1_share1_reg , x0x1x2x3_subscript1_share1_reg , x0x1x2x5_subscript1_share1_reg , x0x1x2x6_subscript1_share1_reg , x0x1x2x7_subscript1_share1_reg , x0x1x4x5_subscript1_share1_reg , x0x1x4x7_subscript1_share1_reg , x0x2x3x5_subscript1_share1_reg , x0x2x3x7_subscript1_share1_reg , x0x2x4x5_subscript1_share1_reg , x0x2x4x7_subscript1_share1_reg , x0x2x5x6_subscript1_share1_reg , x0x2x5x7_subscript1_share1_reg , x0x3x4x6_subscript1_share1_reg , x0x3x5x6_subscript1_share1_reg , x0x4x5x6_subscript1_share1_reg , x0x4x5x7_subscript1_share1_reg , x0x4x6x7_subscript1_share1_reg , x1x2x3x5_subscript1_share1_reg , x1x2x3x6_subscript1_share1_reg , x1x2x3x7_subscript1_share1_reg , x1x2x4x6_subscript1_share1_reg , x1x2x4x7_subscript1_share1_reg , x1x2x6x7_subscript1_share1_reg , x1x3x4x6_subscript1_share1_reg , x1x3x6x7_subscript1_share1_reg , x1x4x5x6_subscript1_share1_reg , x1x4x5x7_subscript1_share1_reg , x1x5x6x7_subscript1_share1_reg , x2x3x5x7_subscript1_share1_reg , x2x3x6x7_subscript1_share1_reg , x2x4x5x6_subscript1_share1_reg , x2x4x5x7_subscript1_share1_reg , x3x5x6x7_subscript1_share1_reg , x0x1x3x4_subscript1_share1_reg , x0x1x3x6_subscript1_share1_reg , x0x1x5x6_subscript1_share1_reg , x0x2x3x6_subscript1_share1_reg , x0x3x4x5_subscript1_share1_reg , x1x2x5x6_subscript1_share1_reg , x1x2x5x7_subscript1_share1_reg , x1x3x4x5_subscript1_share1_reg , x1x3x4x7_subscript1_share1_reg , x1x3x5x6_subscript1_share1_reg , x1x3x5x7_subscript1_share1_reg , x1x4x6x7_subscript1_share1_reg , x2x3x4x5_subscript1_share1_reg , x2x3x4x7_subscript1_share1_reg , x2x4x6x7_subscript1_share1_reg , x3x4x5x6_subscript1_share1_reg , x3x4x5x7_subscript1_share1_reg , x3x4x6x7_subscript1_share1_reg , x0x1x3x5_subscript1_share1_reg , x0x1x4x6_subscript1_share1_reg , x0x2x3x4_subscript1_share1_reg , x0x2x4x6_subscript1_share1_reg , x0x3x4x7_subscript1_share1_reg , x0x3x5x7_subscript1_share1_reg , x1x2x3x4_subscript1_share1_reg , x2x3x4x6_subscript1_share1_reg , x2x3x5x6_subscript1_share1_reg , x2x5x6x7_subscript1_share1_reg , x4x5x6x7_subscript1_share1_reg , x0x1x2x4_subscript1_share1_reg , x0x1x6x7_subscript1_share1_reg , x0x2x6x7_subscript1_share1_reg , x0x3x6x7_subscript1_share1_reg , x0x5x6x7_subscript1_share1_reg , x1x2x4x5_subscript1_share1_reg , x0x1x3x7_subscript1_share1_reg , x0x1x5x7_subscript1_share1_reg , x0x1x2x3x4_subscript1_share1_reg , x0x1x2x3x6_subscript1_share1_reg , x0x1x2x3x7_subscript1_share1_reg , x0x1x2x4x5_subscript1_share1_reg , x0x1x2x4x7_subscript1_share1_reg , x0x1x2x5x7_subscript1_share1_reg , x0x1x2x6x7_subscript1_share1_reg , x0x1x3x4x6_subscript1_share1_reg , x0x1x3x5x6_subscript1_share1_reg , x0x1x3x5x7_subscript1_share1_reg , x0x1x3x6x7_subscript1_share1_reg , x0x1x4x5x6_subscript1_share1_reg , x0x1x5x6x7_subscript1_share1_reg , x0x2x3x4x5_subscript1_share1_reg , x0x2x3x4x6_subscript1_share1_reg , x0x2x4x5x7_subscript1_share1_reg , x0x2x4x6x7_subscript1_share1_reg , x0x3x4x5x6_subscript1_share1_reg , x0x3x4x5x7_subscript1_share1_reg , x0x3x4x6x7_subscript1_share1_reg , x0x3x5x6x7_subscript1_share1_reg , x1x2x3x5x6_subscript1_share1_reg , x1x2x3x5x7_subscript1_share1_reg , x1x2x4x5x6_subscript1_share1_reg , x1x2x4x6x7_subscript1_share1_reg , x1x2x5x6x7_subscript1_share1_reg , x1x3x4x5x7_subscript1_share1_reg , x2x3x4x5x6_subscript1_share1_reg , x2x3x4x5x7_subscript1_share1_reg , x2x4x5x6x7_subscript1_share1_reg , x0x1x2x4x6_subscript1_share1_reg , x0x1x3x4x7_subscript1_share1_reg , x0x2x3x4x7_subscript1_share1_reg , x0x2x3x5x7_subscript1_share1_reg , x0x2x3x6x7_subscript1_share1_reg , x0x2x4x5x6_subscript1_share1_reg , x0x2x5x6x7_subscript1_share1_reg , x0x4x5x6x7_subscript1_share1_reg , x1x2x3x4x6_subscript1_share1_reg , x1x3x4x5x6_subscript1_share1_reg , x2x3x4x6x7_subscript1_share1_reg , x0x1x2x3x5_subscript1_share1_reg , x0x1x4x6x7_subscript1_share1_reg , x1x2x3x4x5_subscript1_share1_reg , x1x2x3x6x7_subscript1_share1_reg , x1x2x4x5x7_subscript1_share1_reg , x1x3x4x6x7_subscript1_share1_reg , x1x3x5x6x7_subscript1_share1_reg , x1x4x5x6x7_subscript1_share1_reg , x2x3x5x6x7_subscript1_share1_reg , x3x4x5x6x7_subscript1_share1_reg , x0x1x2x5x6_subscript1_share1_reg , x0x1x3x4x5_subscript1_share1_reg , x0x1x4x5x7_subscript1_share1_reg , x0x2x3x5x6_subscript1_share1_reg , x1x2x3x4x7_subscript1_share1_reg , x0x1x2x3x4x6_subscript1_share1_reg , x0x1x2x3x4x7_subscript1_share1_reg , x0x1x2x3x5x7_subscript1_share1_reg , x0x1x2x3x6x7_subscript1_share1_reg , x0x1x2x4x5x7_subscript1_share1_reg , x0x1x2x5x6x7_subscript1_share1_reg , x0x1x3x4x6x7_subscript1_share1_reg , x0x1x4x5x6x7_subscript1_share1_reg , x0x2x3x4x5x6_subscript1_share1_reg , x0x2x3x4x5x7_subscript1_share1_reg , x0x2x3x5x6x7_subscript1_share1_reg , x1x2x3x4x6x7_subscript1_share1_reg , x1x2x4x5x6x7_subscript1_share1_reg , x1x3x4x5x6x7_subscript1_share1_reg , x2x3x4x5x6x7_subscript1_share1_reg , x0x1x2x3x5x6_subscript1_share1_reg , x0x1x2x4x6x7_subscript1_share1_reg , x0x1x3x4x5x6_subscript1_share1_reg , x0x2x3x4x6x7_subscript1_share1_reg , x1x2x3x4x5x6_subscript1_share1_reg , x1x2x3x5x6x7_subscript1_share1_reg , x0x1x2x3x4x5_subscript1_share1_reg , x0x1x2x4x5x6_subscript1_share1_reg , x0x1x3x4x5x7_subscript1_share1_reg , x0x1x3x5x6x7_subscript1_share1_reg , x0x2x4x5x6x7_subscript1_share1_reg , x1x2x3x4x5x7_subscript1_share1_reg , x0x3x4x5x6x7_subscript1_share1_reg , x0x1x2x3x4x6x7_subscript1_share1_reg , x0x1x2x4x5x6x7_subscript1_share1_reg , x0x2x3x4x5x6x7_subscript1_share1_reg , x0x1x2x3x5x6x7_subscript1_share1_reg , x0x1x3x4x5x6x7_subscript1_share1_reg , x1x2x3x4x5x6x7_subscript1_share1_reg , x0x1x2x3x4x5x6_subscript1_share1_reg , x0x1x2x3x4x5x7_subscript1_share1_reg , 
    x0_pipelined2_share3_reg ,x1_pipelined2_share3_reg ,x2_pipelined2_share3_reg ,x3_pipelined2_share3_reg ,x4_pipelined2_share3_reg ,x5_pipelined2_share3_reg ,x6_pipelined2_share3_reg ,x7_pipelined2_share3_reg ,
    sbox_out1_share1, sbox_out2_share1, sbox_out3_share1, sbox_out4_share1, sbox_out5_share1, sbox_out6_share1, sbox_out7_share1, sbox_out8_share1 
);

combi_logic_cycle3_output_share2 inst_cycle3_share2 (
    x0_subscript1_share2_reg , x2_subscript1_share2_reg , x3_subscript1_share2_reg , x4_subscript1_share2_reg , x6_subscript1_share2_reg , x7_subscript1_share2_reg , x1_subscript1_share2_reg , x5_subscript1_share2_reg , x0x1_subscript1_share2_reg , x0x4_subscript1_share2_reg , x0x5_subscript1_share2_reg , x0x6_subscript1_share2_reg , x1x2_subscript1_share2_reg , x1x3_subscript1_share2_reg , x1x4_subscript1_share2_reg , x1x6_subscript1_share2_reg , x2x3_subscript1_share2_reg , x2x4_subscript1_share2_reg , x2x6_subscript1_share2_reg , x2x7_subscript1_share2_reg , x4x6_subscript1_share2_reg , x5x6_subscript1_share2_reg , x5x7_subscript1_share2_reg , x6x7_subscript1_share2_reg , x0x2_subscript1_share2_reg , x0x3_subscript1_share2_reg , x0x7_subscript1_share2_reg , x1x7_subscript1_share2_reg , x3x7_subscript1_share2_reg , x4x5_subscript1_share2_reg , x3x4_subscript1_share2_reg , x4x7_subscript1_share2_reg , x3x6_subscript1_share2_reg , x1x5_subscript1_share2_reg , x2x5_subscript1_share2_reg , x3x5_subscript1_share2_reg , x0x1x4_subscript1_share2_reg , x0x1x6_subscript1_share2_reg , x0x1x7_subscript1_share2_reg , x0x2x4_subscript1_share2_reg , x0x2x5_subscript1_share2_reg , x0x2x6_subscript1_share2_reg , x0x2x7_subscript1_share2_reg , x0x3x4_subscript1_share2_reg , x0x3x5_subscript1_share2_reg , x0x3x6_subscript1_share2_reg , x0x4x6_subscript1_share2_reg , x0x4x7_subscript1_share2_reg , x1x2x3_subscript1_share2_reg , x1x2x4_subscript1_share2_reg , x1x2x6_subscript1_share2_reg , x1x3x4_subscript1_share2_reg , x1x3x7_subscript1_share2_reg , x1x4x6_subscript1_share2_reg , x1x5x6_subscript1_share2_reg , x2x3x5_subscript1_share2_reg , x2x3x7_subscript1_share2_reg , x2x4x7_subscript1_share2_reg , x2x5x6_subscript1_share2_reg , x2x5x7_subscript1_share2_reg , x2x6x7_subscript1_share2_reg , x3x4x7_subscript1_share2_reg , x3x5x7_subscript1_share2_reg , x3x6x7_subscript1_share2_reg , x4x5x6_subscript1_share2_reg , x5x6x7_subscript1_share2_reg , x0x1x3_subscript1_share2_reg , x0x2x3_subscript1_share2_reg , x0x4x5_subscript1_share2_reg , x0x5x7_subscript1_share2_reg , x0x6x7_subscript1_share2_reg , x1x3x5_subscript1_share2_reg , x1x3x6_subscript1_share2_reg , x1x4x7_subscript1_share2_reg , x2x3x4_subscript1_share2_reg , x2x3x6_subscript1_share2_reg , x3x4x6_subscript1_share2_reg , x3x5x6_subscript1_share2_reg , x0x1x5_subscript1_share2_reg , x0x3x7_subscript1_share2_reg , x1x2x5_subscript1_share2_reg , x1x2x7_subscript1_share2_reg , x1x4x5_subscript1_share2_reg , x1x5x7_subscript1_share2_reg , x2x4x5_subscript1_share2_reg , x3x4x5_subscript1_share2_reg , x4x6x7_subscript1_share2_reg , x1x6x7_subscript1_share2_reg , x4x5x7_subscript1_share2_reg , x0x1x2_subscript1_share2_reg , x0x5x6_subscript1_share2_reg , x2x4x6_subscript1_share2_reg , x0x1x2x3_subscript1_share2_reg , x0x1x2x5_subscript1_share2_reg , x0x1x2x6_subscript1_share2_reg , x0x1x2x7_subscript1_share2_reg , x0x1x4x5_subscript1_share2_reg , x0x1x4x7_subscript1_share2_reg , x0x2x3x5_subscript1_share2_reg , x0x2x3x7_subscript1_share2_reg , x0x2x4x5_subscript1_share2_reg , x0x2x4x7_subscript1_share2_reg , x0x2x5x6_subscript1_share2_reg , x0x2x5x7_subscript1_share2_reg , x0x3x4x6_subscript1_share2_reg , x0x3x5x6_subscript1_share2_reg , x0x4x5x6_subscript1_share2_reg , x0x4x5x7_subscript1_share2_reg , x0x4x6x7_subscript1_share2_reg , x1x2x3x5_subscript1_share2_reg , x1x2x3x6_subscript1_share2_reg , x1x2x3x7_subscript1_share2_reg , x1x2x4x6_subscript1_share2_reg , x1x2x4x7_subscript1_share2_reg , x1x2x6x7_subscript1_share2_reg , x1x3x4x6_subscript1_share2_reg , x1x3x6x7_subscript1_share2_reg , x1x4x5x6_subscript1_share2_reg , x1x4x5x7_subscript1_share2_reg , x1x5x6x7_subscript1_share2_reg , x2x3x5x7_subscript1_share2_reg , x2x3x6x7_subscript1_share2_reg , x2x4x5x6_subscript1_share2_reg , x2x4x5x7_subscript1_share2_reg , x3x5x6x7_subscript1_share2_reg , x0x1x3x4_subscript1_share2_reg , x0x1x3x6_subscript1_share2_reg , x0x1x5x6_subscript1_share2_reg , x0x2x3x6_subscript1_share2_reg , x0x3x4x5_subscript1_share2_reg , x1x2x5x6_subscript1_share2_reg , x1x2x5x7_subscript1_share2_reg , x1x3x4x5_subscript1_share2_reg , x1x3x4x7_subscript1_share2_reg , x1x3x5x6_subscript1_share2_reg , x1x3x5x7_subscript1_share2_reg , x1x4x6x7_subscript1_share2_reg , x2x3x4x5_subscript1_share2_reg , x2x3x4x7_subscript1_share2_reg , x2x4x6x7_subscript1_share2_reg , x3x4x5x6_subscript1_share2_reg , x3x4x5x7_subscript1_share2_reg , x3x4x6x7_subscript1_share2_reg , x0x1x3x5_subscript1_share2_reg , x0x1x4x6_subscript1_share2_reg , x0x2x3x4_subscript1_share2_reg , x0x2x4x6_subscript1_share2_reg , x0x3x4x7_subscript1_share2_reg , x0x3x5x7_subscript1_share2_reg , x1x2x3x4_subscript1_share2_reg , x2x3x4x6_subscript1_share2_reg , x2x3x5x6_subscript1_share2_reg , x2x5x6x7_subscript1_share2_reg , x4x5x6x7_subscript1_share2_reg , x0x1x2x4_subscript1_share2_reg , x0x1x6x7_subscript1_share2_reg , x0x2x6x7_subscript1_share2_reg , x0x3x6x7_subscript1_share2_reg , x0x5x6x7_subscript1_share2_reg , x1x2x4x5_subscript1_share2_reg , x0x1x3x7_subscript1_share2_reg , x0x1x5x7_subscript1_share2_reg , x0x1x2x3x4_subscript1_share2_reg , x0x1x2x3x6_subscript1_share2_reg , x0x1x2x3x7_subscript1_share2_reg , x0x1x2x4x5_subscript1_share2_reg , x0x1x2x4x7_subscript1_share2_reg , x0x1x2x5x7_subscript1_share2_reg , x0x1x2x6x7_subscript1_share2_reg , x0x1x3x4x6_subscript1_share2_reg , x0x1x3x5x6_subscript1_share2_reg , x0x1x3x5x7_subscript1_share2_reg , x0x1x3x6x7_subscript1_share2_reg , x0x1x4x5x6_subscript1_share2_reg , x0x1x5x6x7_subscript1_share2_reg , x0x2x3x4x5_subscript1_share2_reg , x0x2x3x4x6_subscript1_share2_reg , x0x2x4x5x7_subscript1_share2_reg , x0x2x4x6x7_subscript1_share2_reg , x0x3x4x5x6_subscript1_share2_reg , x0x3x4x5x7_subscript1_share2_reg , x0x3x4x6x7_subscript1_share2_reg , x0x3x5x6x7_subscript1_share2_reg , x1x2x3x5x6_subscript1_share2_reg , x1x2x3x5x7_subscript1_share2_reg , x1x2x4x5x6_subscript1_share2_reg , x1x2x4x6x7_subscript1_share2_reg , x1x2x5x6x7_subscript1_share2_reg , x1x3x4x5x7_subscript1_share2_reg , x2x3x4x5x6_subscript1_share2_reg , x2x3x4x5x7_subscript1_share2_reg , x2x4x5x6x7_subscript1_share2_reg , x0x1x2x4x6_subscript1_share2_reg , x0x1x3x4x7_subscript1_share2_reg , x0x2x3x4x7_subscript1_share2_reg , x0x2x3x5x7_subscript1_share2_reg , x0x2x3x6x7_subscript1_share2_reg , x0x2x4x5x6_subscript1_share2_reg , x0x2x5x6x7_subscript1_share2_reg , x0x4x5x6x7_subscript1_share2_reg , x1x2x3x4x6_subscript1_share2_reg , x1x3x4x5x6_subscript1_share2_reg , x2x3x4x6x7_subscript1_share2_reg , x0x1x2x3x5_subscript1_share2_reg , x0x1x4x6x7_subscript1_share2_reg , x1x2x3x4x5_subscript1_share2_reg , x1x2x3x6x7_subscript1_share2_reg , x1x2x4x5x7_subscript1_share2_reg , x1x3x4x6x7_subscript1_share2_reg , x1x3x5x6x7_subscript1_share2_reg , x1x4x5x6x7_subscript1_share2_reg , x2x3x5x6x7_subscript1_share2_reg , x3x4x5x6x7_subscript1_share2_reg , x0x1x2x5x6_subscript1_share2_reg , x0x1x3x4x5_subscript1_share2_reg , x0x1x4x5x7_subscript1_share2_reg , x0x2x3x5x6_subscript1_share2_reg , x1x2x3x4x7_subscript1_share2_reg , x0x1x2x3x4x6_subscript1_share2_reg , x0x1x2x3x4x7_subscript1_share2_reg , x0x1x2x3x5x7_subscript1_share2_reg , x0x1x2x3x6x7_subscript1_share2_reg , x0x1x2x4x5x7_subscript1_share2_reg , x0x1x2x5x6x7_subscript1_share2_reg , x0x1x3x4x6x7_subscript1_share2_reg , x0x1x4x5x6x7_subscript1_share2_reg , x0x2x3x4x5x6_subscript1_share2_reg , x0x2x3x4x5x7_subscript1_share2_reg , x0x2x3x5x6x7_subscript1_share2_reg , x1x2x3x4x6x7_subscript1_share2_reg , x1x2x4x5x6x7_subscript1_share2_reg , x1x3x4x5x6x7_subscript1_share2_reg , x2x3x4x5x6x7_subscript1_share2_reg , x0x1x2x3x5x6_subscript1_share2_reg , x0x1x2x4x6x7_subscript1_share2_reg , x0x1x3x4x5x6_subscript1_share2_reg , x0x2x3x4x6x7_subscript1_share2_reg , x1x2x3x4x5x6_subscript1_share2_reg , x1x2x3x5x6x7_subscript1_share2_reg , x0x1x2x3x4x5_subscript1_share2_reg , x0x1x2x4x5x6_subscript1_share2_reg , x0x1x3x4x5x7_subscript1_share2_reg , x0x1x3x5x6x7_subscript1_share2_reg , x0x2x4x5x6x7_subscript1_share2_reg , x1x2x3x4x5x7_subscript1_share2_reg , x0x3x4x5x6x7_subscript1_share2_reg , x0x1x2x3x4x6x7_subscript1_share2_reg , x0x1x2x4x5x6x7_subscript1_share2_reg , x0x2x3x4x5x6x7_subscript1_share2_reg , x0x1x2x3x5x6x7_subscript1_share2_reg , x0x1x3x4x5x6x7_subscript1_share2_reg , x1x2x3x4x5x6x7_subscript1_share2_reg , x0x1x2x3x4x5x6_subscript1_share2_reg , x0x1x2x3x4x5x7_subscript1_share2_reg , 
    x0_pipelined2_share3_reg ,x1_pipelined2_share3_reg ,x2_pipelined2_share3_reg ,x3_pipelined2_share3_reg ,x4_pipelined2_share3_reg ,x5_pipelined2_share3_reg ,x6_pipelined2_share3_reg ,x7_pipelined2_share3_reg ,
    sbox_out1_share2, sbox_out2_share2, sbox_out3_share2, sbox_out4_share2, sbox_out5_share2, sbox_out6_share2, sbox_out7_share2, sbox_out8_share2 
);

combi_logic_cycle3_output_share3 inst_cycle3_share3 (
    x0_subscript1_share3_reg , x2_subscript1_share3_reg , x3_subscript1_share3_reg , x4_subscript1_share3_reg , x6_subscript1_share3_reg , x7_subscript1_share3_reg , x1_subscript1_share3_reg , x5_subscript1_share3_reg , x0x1_subscript1_share3_reg , x0x4_subscript1_share3_reg , x0x5_subscript1_share3_reg , x0x6_subscript1_share3_reg , x1x2_subscript1_share3_reg , x1x3_subscript1_share3_reg , x1x4_subscript1_share3_reg , x1x6_subscript1_share3_reg , x2x3_subscript1_share3_reg , x2x4_subscript1_share3_reg , x2x6_subscript1_share3_reg , x2x7_subscript1_share3_reg , x4x6_subscript1_share3_reg , x5x6_subscript1_share3_reg , x5x7_subscript1_share3_reg , x6x7_subscript1_share3_reg , x0x2_subscript1_share3_reg , x0x3_subscript1_share3_reg , x0x7_subscript1_share3_reg , x1x7_subscript1_share3_reg , x3x7_subscript1_share3_reg , x4x5_subscript1_share3_reg , x3x4_subscript1_share3_reg , x4x7_subscript1_share3_reg , x3x6_subscript1_share3_reg , x1x5_subscript1_share3_reg , x2x5_subscript1_share3_reg , x3x5_subscript1_share3_reg , x0x1x4_subscript1_share3_reg , x0x1x6_subscript1_share3_reg , x0x1x7_subscript1_share3_reg , x0x2x4_subscript1_share3_reg , x0x2x5_subscript1_share3_reg , x0x2x6_subscript1_share3_reg , x0x2x7_subscript1_share3_reg , x0x3x4_subscript1_share3_reg , x0x3x5_subscript1_share3_reg , x0x3x6_subscript1_share3_reg , x0x4x6_subscript1_share3_reg , x0x4x7_subscript1_share3_reg , x1x2x3_subscript1_share3_reg , x1x2x4_subscript1_share3_reg , x1x2x6_subscript1_share3_reg , x1x3x4_subscript1_share3_reg , x1x3x7_subscript1_share3_reg , x1x4x6_subscript1_share3_reg , x1x5x6_subscript1_share3_reg , x2x3x5_subscript1_share3_reg , x2x3x7_subscript1_share3_reg , x2x4x7_subscript1_share3_reg , x2x5x6_subscript1_share3_reg , x2x5x7_subscript1_share3_reg , x2x6x7_subscript1_share3_reg , x3x4x7_subscript1_share3_reg , x3x5x7_subscript1_share3_reg , x3x6x7_subscript1_share3_reg , x4x5x6_subscript1_share3_reg , x5x6x7_subscript1_share3_reg , x0x1x3_subscript1_share3_reg , x0x2x3_subscript1_share3_reg , x0x4x5_subscript1_share3_reg , x0x5x7_subscript1_share3_reg , x0x6x7_subscript1_share3_reg , x1x3x5_subscript1_share3_reg , x1x3x6_subscript1_share3_reg , x1x4x7_subscript1_share3_reg , x2x3x4_subscript1_share3_reg , x2x3x6_subscript1_share3_reg , x3x4x6_subscript1_share3_reg , x3x5x6_subscript1_share3_reg , x0x1x5_subscript1_share3_reg , x0x3x7_subscript1_share3_reg , x1x2x5_subscript1_share3_reg , x1x2x7_subscript1_share3_reg , x1x4x5_subscript1_share3_reg , x1x5x7_subscript1_share3_reg , x2x4x5_subscript1_share3_reg , x3x4x5_subscript1_share3_reg , x4x6x7_subscript1_share3_reg , x1x6x7_subscript1_share3_reg , x4x5x7_subscript1_share3_reg , x0x1x2_subscript1_share3_reg , x0x5x6_subscript1_share3_reg , x2x4x6_subscript1_share3_reg , x0x1x2x3_subscript1_share3_reg , x0x1x2x5_subscript1_share3_reg , x0x1x2x6_subscript1_share3_reg , x0x1x2x7_subscript1_share3_reg , x0x1x4x5_subscript1_share3_reg , x0x1x4x7_subscript1_share3_reg , x0x2x3x5_subscript1_share3_reg , x0x2x3x7_subscript1_share3_reg , x0x2x4x5_subscript1_share3_reg , x0x2x4x7_subscript1_share3_reg , x0x2x5x6_subscript1_share3_reg , x0x2x5x7_subscript1_share3_reg , x0x3x4x6_subscript1_share3_reg , x0x3x5x6_subscript1_share3_reg , x0x4x5x6_subscript1_share3_reg , x0x4x5x7_subscript1_share3_reg , x0x4x6x7_subscript1_share3_reg , x1x2x3x5_subscript1_share3_reg , x1x2x3x6_subscript1_share3_reg , x1x2x3x7_subscript1_share3_reg , x1x2x4x6_subscript1_share3_reg , x1x2x4x7_subscript1_share3_reg , x1x2x6x7_subscript1_share3_reg , x1x3x4x6_subscript1_share3_reg , x1x3x6x7_subscript1_share3_reg , x1x4x5x6_subscript1_share3_reg , x1x4x5x7_subscript1_share3_reg , x1x5x6x7_subscript1_share3_reg , x2x3x5x7_subscript1_share3_reg , x2x3x6x7_subscript1_share3_reg , x2x4x5x6_subscript1_share3_reg , x2x4x5x7_subscript1_share3_reg , x3x5x6x7_subscript1_share3_reg , x0x1x3x4_subscript1_share3_reg , x0x1x3x6_subscript1_share3_reg , x0x1x5x6_subscript1_share3_reg , x0x2x3x6_subscript1_share3_reg , x0x3x4x5_subscript1_share3_reg , x1x2x5x6_subscript1_share3_reg , x1x2x5x7_subscript1_share3_reg , x1x3x4x5_subscript1_share3_reg , x1x3x4x7_subscript1_share3_reg , x1x3x5x6_subscript1_share3_reg , x1x3x5x7_subscript1_share3_reg , x1x4x6x7_subscript1_share3_reg , x2x3x4x5_subscript1_share3_reg , x2x3x4x7_subscript1_share3_reg , x2x4x6x7_subscript1_share3_reg , x3x4x5x6_subscript1_share3_reg , x3x4x5x7_subscript1_share3_reg , x3x4x6x7_subscript1_share3_reg , x0x1x3x5_subscript1_share3_reg , x0x1x4x6_subscript1_share3_reg , x0x2x3x4_subscript1_share3_reg , x0x2x4x6_subscript1_share3_reg , x0x3x4x7_subscript1_share3_reg , x0x3x5x7_subscript1_share3_reg , x1x2x3x4_subscript1_share3_reg , x2x3x4x6_subscript1_share3_reg , x2x3x5x6_subscript1_share3_reg , x2x5x6x7_subscript1_share3_reg , x4x5x6x7_subscript1_share3_reg , x0x1x2x4_subscript1_share3_reg , x0x1x6x7_subscript1_share3_reg , x0x2x6x7_subscript1_share3_reg , x0x3x6x7_subscript1_share3_reg , x0x5x6x7_subscript1_share3_reg , x1x2x4x5_subscript1_share3_reg , x0x1x3x7_subscript1_share3_reg , x0x1x5x7_subscript1_share3_reg , x0x1x2x3x4_subscript1_share3_reg , x0x1x2x3x6_subscript1_share3_reg , x0x1x2x3x7_subscript1_share3_reg , x0x1x2x4x5_subscript1_share3_reg , x0x1x2x4x7_subscript1_share3_reg , x0x1x2x5x7_subscript1_share3_reg , x0x1x2x6x7_subscript1_share3_reg , x0x1x3x4x6_subscript1_share3_reg , x0x1x3x5x6_subscript1_share3_reg , x0x1x3x5x7_subscript1_share3_reg , x0x1x3x6x7_subscript1_share3_reg , x0x1x4x5x6_subscript1_share3_reg , x0x1x5x6x7_subscript1_share3_reg , x0x2x3x4x5_subscript1_share3_reg , x0x2x3x4x6_subscript1_share3_reg , x0x2x4x5x7_subscript1_share3_reg , x0x2x4x6x7_subscript1_share3_reg , x0x3x4x5x6_subscript1_share3_reg , x0x3x4x5x7_subscript1_share3_reg , x0x3x4x6x7_subscript1_share3_reg , x0x3x5x6x7_subscript1_share3_reg , x1x2x3x5x6_subscript1_share3_reg , x1x2x3x5x7_subscript1_share3_reg , x1x2x4x5x6_subscript1_share3_reg , x1x2x4x6x7_subscript1_share3_reg , x1x2x5x6x7_subscript1_share3_reg , x1x3x4x5x7_subscript1_share3_reg , x2x3x4x5x6_subscript1_share3_reg , x2x3x4x5x7_subscript1_share3_reg , x2x4x5x6x7_subscript1_share3_reg , x0x1x2x4x6_subscript1_share3_reg , x0x1x3x4x7_subscript1_share3_reg , x0x2x3x4x7_subscript1_share3_reg , x0x2x3x5x7_subscript1_share3_reg , x0x2x3x6x7_subscript1_share3_reg , x0x2x4x5x6_subscript1_share3_reg , x0x2x5x6x7_subscript1_share3_reg , x0x4x5x6x7_subscript1_share3_reg , x1x2x3x4x6_subscript1_share3_reg , x1x3x4x5x6_subscript1_share3_reg , x2x3x4x6x7_subscript1_share3_reg , x0x1x2x3x5_subscript1_share3_reg , x0x1x4x6x7_subscript1_share3_reg , x1x2x3x4x5_subscript1_share3_reg , x1x2x3x6x7_subscript1_share3_reg , x1x2x4x5x7_subscript1_share3_reg , x1x3x4x6x7_subscript1_share3_reg , x1x3x5x6x7_subscript1_share3_reg , x1x4x5x6x7_subscript1_share3_reg , x2x3x5x6x7_subscript1_share3_reg , x3x4x5x6x7_subscript1_share3_reg , x0x1x2x5x6_subscript1_share3_reg , x0x1x3x4x5_subscript1_share3_reg , x0x1x4x5x7_subscript1_share3_reg , x0x2x3x5x6_subscript1_share3_reg , x1x2x3x4x7_subscript1_share3_reg , x0x1x2x3x4x6_subscript1_share3_reg , x0x1x2x3x4x7_subscript1_share3_reg , x0x1x2x3x5x7_subscript1_share3_reg , x0x1x2x3x6x7_subscript1_share3_reg , x0x1x2x4x5x7_subscript1_share3_reg , x0x1x2x5x6x7_subscript1_share3_reg , x0x1x3x4x6x7_subscript1_share3_reg , x0x1x4x5x6x7_subscript1_share3_reg , x0x2x3x4x5x6_subscript1_share3_reg , x0x2x3x4x5x7_subscript1_share3_reg , x0x2x3x5x6x7_subscript1_share3_reg , x1x2x3x4x6x7_subscript1_share3_reg , x1x2x4x5x6x7_subscript1_share3_reg , x1x3x4x5x6x7_subscript1_share3_reg , x2x3x4x5x6x7_subscript1_share3_reg , x0x1x2x3x5x6_subscript1_share3_reg , x0x1x2x4x6x7_subscript1_share3_reg , x0x1x3x4x5x6_subscript1_share3_reg , x0x2x3x4x6x7_subscript1_share3_reg , x1x2x3x4x5x6_subscript1_share3_reg , x1x2x3x5x6x7_subscript1_share3_reg , x0x1x2x3x4x5_subscript1_share3_reg , x0x1x2x4x5x6_subscript1_share3_reg , x0x1x3x4x5x7_subscript1_share3_reg , x0x1x3x5x6x7_subscript1_share3_reg , x0x2x4x5x6x7_subscript1_share3_reg , x1x2x3x4x5x7_subscript1_share3_reg , x0x3x4x5x6x7_subscript1_share3_reg , x0x1x2x3x4x6x7_subscript1_share3_reg , x0x1x2x4x5x6x7_subscript1_share3_reg , x0x2x3x4x5x6x7_subscript1_share3_reg , x0x1x2x3x5x6x7_subscript1_share3_reg , x0x1x3x4x5x6x7_subscript1_share3_reg , x1x2x3x4x5x6x7_subscript1_share3_reg , x0x1x2x3x4x5x6_subscript1_share3_reg , x0x1x2x3x4x5x7_subscript1_share3_reg , 
    x0_pipelined2_share3_reg ,x1_pipelined2_share3_reg ,x2_pipelined2_share3_reg ,x3_pipelined2_share3_reg ,x4_pipelined2_share3_reg ,x5_pipelined2_share3_reg ,x6_pipelined2_share3_reg ,x7_pipelined2_share3_reg ,
    sbox_out1_share3, sbox_out2_share3, sbox_out3_share3, sbox_out4_share3, sbox_out5_share3, sbox_out6_share3, sbox_out7_share3, sbox_out8_share3 
);

assign output_share1 = {sbox_out8_share1, sbox_out7_share1, sbox_out6_share1, sbox_out5_share1, sbox_out4_share1, sbox_out3_share1, sbox_out2_share1, sbox_out1_share1} ;
assign output_share2 = {sbox_out8_share2, sbox_out7_share2, sbox_out6_share2, sbox_out5_share2, sbox_out4_share2, sbox_out3_share2, sbox_out2_share2, sbox_out1_share2} ;
assign output_share3 = {sbox_out8_share3, sbox_out7_share3, sbox_out6_share3, sbox_out5_share3, sbox_out4_share3, sbox_out3_share3, sbox_out2_share3, sbox_out1_share3} ;


endmodule