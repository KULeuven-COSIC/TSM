`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 22:00:00 02/22/2025
// Design Name: Register Array for One Share
// Module Name: register_array_AES_oneshare
// Project Name: AES Masked S-Box
// Description: Stores 254 input signals using registers and outputs stored values for exactly one share.
// Dependencies: None
//
// Revision:
// Revision 0.01 - Initial version
//
//////////////////////////////////////////////////////////////////////////////////


module register_array_AES_oneshare(
clk,
in1 , in2 , in3 , in4 , in5 , in6 , in7 , in8 , in9 , in10 , in11 , in12 , in13 , in14 , in15 , in16 , in17 , in18 , in19 , in20 , in21 , in22 , in23 , in24 , in25 , in26 , in27 , in28 , in29 , in30 , in31 , in32 , in33 , in34 , in35 , in36 , in37 , in38 , in39 , in40 , in41 , in42 , in43 , in44 , in45 , in46 , in47 , in48 , in49 , in50 , in51 , in52 , in53 , in54 , in55 , in56 , in57 , in58 , in59 , in60 , in61 , in62 , in63 , in64 , in65 , in66 , in67 , in68 , in69 , in70 , in71 , in72 , in73 , in74 , in75 , in76 , in77 , in78 , in79 , in80 , in81 , in82 , in83 , in84 , in85 , in86 , in87 , in88 , in89 , in90 , in91 , in92 , in93 , in94 , in95 , in96 , in97 , in98 , in99 , in100 , in101 , in102 , in103 , in104 , in105 , in106 , in107 , in108 , in109 , in110 , in111 , in112 , in113 , in114 , in115 , in116 , in117 , in118 , in119 , in120 , in121 , in122 , in123 , in124 , in125 , in126 , in127 , in128 , in129 , in130 , in131 , in132 , in133 , in134 , in135 , in136 , in137 , in138 , in139 , in140 , in141 , in142 , in143 , in144 , in145 , in146 , in147 , in148 , in149 , in150 , in151 , in152 , in153 , in154 , in155 , in156 , in157 , in158 , in159 , in160 , in161 , in162 , in163 , in164 , in165 , in166 , in167 , in168 , in169 , in170 , in171 , in172 , in173 , in174 , in175 , in176 , in177 , in178 , in179 , in180 , in181 , in182 , in183 , in184 , in185 , in186 , in187 , in188 , in189 , in190 , in191 , in192 , in193 , in194 , in195 , in196 , in197 , in198 , in199 , in200 , in201 , in202 , in203 , in204 , in205 , in206 , in207 , in208 , in209 , in210 , in211 , in212 , in213 , in214 , in215 , in216 , in217 , in218 , in219 , in220 , in221 , in222 , in223 , in224 , in225 , in226 , in227 , in228 , in229 , in230 , in231 , in232 , in233 , in234 , in235 , in236 , in237 , in238 , in239 , in240 , in241 , in242 , in243 , in244 , in245 , in246 , in247 , in248 , in249 , in250 , in251 , in252 , in253 , in254 , 
out1 , out2 , out3 , out4 , out5 , out6 , out7 , out8 , out9 , out10 , out11 , out12 , out13 , out14 , out15 , out16 , out17 , out18 , out19 , out20 , out21 , out22 , out23 , out24 , out25 , out26 , out27 , out28 , out29 , out30 , out31 , out32 , out33 , out34 , out35 , out36 , out37 , out38 , out39 , out40 , out41 , out42 , out43 , out44 , out45 , out46 , out47 , out48 , out49 , out50 , out51 , out52 , out53 , out54 , out55 , out56 , out57 , out58 , out59 , out60 , out61 , out62 , out63 , out64 , out65 , out66 , out67 , out68 , out69 , out70 , out71 , out72 , out73 , out74 , out75 , out76 , out77 , out78 , out79 , out80 , out81 , out82 , out83 , out84 , out85 , out86 , out87 , out88 , out89 , out90 , out91 , out92 , out93 , out94 , out95 , out96 , out97 , out98 , out99 , out100 , out101 , out102 , out103 , out104 , out105 , out106 , out107 , out108 , out109 , out110 , out111 , out112 , out113 , out114 , out115 , out116 , out117 , out118 , out119 , out120 , out121 , out122 , out123 , out124 , out125 , out126 , out127 , out128 , out129 , out130 , out131 , out132 , out133 , out134 , out135 , out136 , out137 , out138 , out139 , out140 , out141 , out142 , out143 , out144 , out145 , out146 , out147 , out148 , out149 , out150 , out151 , out152 , out153 , out154 , out155 , out156 , out157 , out158 , out159 , out160 , out161 , out162 , out163 , out164 , out165 , out166 , out167 , out168 , out169 , out170 , out171 , out172 , out173 , out174 , out175 , out176 , out177 , out178 , out179 , out180 , out181 , out182 , out183 , out184 , out185 , out186 , out187 , out188 , out189 , out190 , out191 , out192 , out193 , out194 , out195 , out196 , out197 , out198 , out199 , out200 , out201 , out202 , out203 , out204 , out205 , out206 , out207 , out208 , out209 , out210 , out211 , out212 , out213 , out214 , out215 , out216 , out217 , out218 , out219 , out220 , out221 , out222 , out223 , out224 , out225 , out226 , out227 , out228 , out229 , out230 , out231 , out232 , out233 , out234 , out235 , out236 , out237 , out238 , out239 , out240 , out241 , out242 , out243 , out244 , out245 , out246 , out247 , out248 , out249 , out250 , out251 , out252 , out253 , out254 
);

input clk ;
input in1 , in2 , in3 , in4 , in5 , in6 , in7 , in8 , in9 , in10 , in11 , in12 , in13 , in14 , in15 , in16 , in17 , in18 , in19 , in20 , in21 , in22 , in23 , in24 , in25 , in26 , in27 , in28 , in29 , in30 , in31 , in32 , in33 , in34 , in35 , in36 , in37 , in38 , in39 , in40 , in41 , in42 , in43 , in44 , in45 , in46 , in47 , in48 , in49 , in50 , in51 , in52 , in53 , in54 , in55 , in56 , in57 , in58 , in59 , in60 , in61 , in62 , in63 , in64 , in65 , in66 , in67 , in68 , in69 , in70 , in71 , in72 , in73 , in74 , in75 , in76 , in77 , in78 , in79 , in80 , in81 , in82 , in83 , in84 , in85 , in86 , in87 , in88 , in89 , in90 , in91 , in92 , in93 , in94 , in95 , in96 , in97 , in98 , in99 , in100 , in101 , in102 , in103 , in104 , in105 , in106 , in107 , in108 , in109 , in110 , in111 , in112 , in113 , in114 , in115 , in116 , in117 , in118 , in119 , in120 , in121 , in122 , in123 , in124 , in125 , in126 , in127 , in128 , in129 , in130 , in131 , in132 , in133 , in134 , in135 , in136 , in137 , in138 , in139 , in140 , in141 , in142 , in143 , in144 , in145 , in146 , in147 , in148 , in149 , in150 , in151 , in152 , in153 , in154 , in155 , in156 , in157 , in158 , in159 , in160 , in161 , in162 , in163 , in164 , in165 , in166 , in167 , in168 , in169 , in170 , in171 , in172 , in173 , in174 , in175 , in176 , in177 , in178 , in179 , in180 , in181 , in182 , in183 , in184 , in185 , in186 , in187 , in188 , in189 , in190 , in191 , in192 , in193 , in194 , in195 , in196 , in197 , in198 , in199 , in200 , in201 , in202 , in203 , in204 , in205 , in206 , in207 , in208 , in209 , in210 , in211 , in212 , in213 , in214 , in215 , in216 , in217 , in218 , in219 , in220 , in221 , in222 , in223 , in224 , in225 , in226 , in227 , in228 , in229 , in230 , in231 , in232 , in233 , in234 , in235 , in236 , in237 , in238 , in239 , in240 , in241 , in242 , in243 , in244 , in245 , in246 , in247 , in248 , in249 , in250 , in251 , in252 , in253 , in254 ;
output out1 , out2 , out3 , out4 , out5 , out6 , out7 , out8 , out9 , out10 , out11 , out12 , out13 , out14 , out15 , out16 , out17 , out18 , out19 , out20 , out21 , out22 , out23 , out24 , out25 , out26 , out27 , out28 , out29 , out30 , out31 , out32 , out33 , out34 , out35 , out36 , out37 , out38 , out39 , out40 , out41 , out42 , out43 , out44 , out45 , out46 , out47 , out48 , out49 , out50 , out51 , out52 , out53 , out54 , out55 , out56 , out57 , out58 , out59 , out60 , out61 , out62 , out63 , out64 , out65 , out66 , out67 , out68 , out69 , out70 , out71 , out72 , out73 , out74 , out75 , out76 , out77 , out78 , out79 , out80 , out81 , out82 , out83 , out84 , out85 , out86 , out87 , out88 , out89 , out90 , out91 , out92 , out93 , out94 , out95 , out96 , out97 , out98 , out99 , out100 , out101 , out102 , out103 , out104 , out105 , out106 , out107 , out108 , out109 , out110 , out111 , out112 , out113 , out114 , out115 , out116 , out117 , out118 , out119 , out120 , out121 , out122 , out123 , out124 , out125 , out126 , out127 , out128 , out129 , out130 , out131 , out132 , out133 , out134 , out135 , out136 , out137 , out138 , out139 , out140 , out141 , out142 , out143 , out144 , out145 , out146 , out147 , out148 , out149 , out150 , out151 , out152 , out153 , out154 , out155 , out156 , out157 , out158 , out159 , out160 , out161 , out162 , out163 , out164 , out165 , out166 , out167 , out168 , out169 , out170 , out171 , out172 , out173 , out174 , out175 , out176 , out177 , out178 , out179 , out180 , out181 , out182 , out183 , out184 , out185 , out186 , out187 , out188 , out189 , out190 , out191 , out192 , out193 , out194 , out195 , out196 , out197 , out198 , out199 , out200 , out201 , out202 , out203 , out204 , out205 , out206 , out207 , out208 , out209 , out210 , out211 , out212 , out213 , out214 , out215 , out216 , out217 , out218 , out219 , out220 , out221 , out222 , out223 , out224 , out225 , out226 , out227 , out228 , out229 , out230 , out231 , out232 , out233 , out234 , out235 , out236 , out237 , out238 , out239 , out240 , out241 , out242 , out243 , out244 , out245 , out246 , out247 , out248 , out249 , out250 , out251 , out252 , out253 , out254  ;

reg  reg_out1 , reg_out2 , reg_out3 , reg_out4 , reg_out5 , reg_out6 , reg_out7 , reg_out8 , reg_out9 , reg_out10 , reg_out11 , reg_out12 , reg_out13 , reg_out14 , reg_out15 , reg_out16 , reg_out17 , reg_out18 , reg_out19 , reg_out20 , reg_out21 , reg_out22 , reg_out23 , reg_out24 , reg_out25 , reg_out26 , reg_out27 , reg_out28 , reg_out29 , reg_out30 , reg_out31 , reg_out32 , reg_out33 , reg_out34 , reg_out35 , reg_out36 , reg_out37 , reg_out38 , reg_out39 , reg_out40 , reg_out41 , reg_out42 , reg_out43 , reg_out44 , reg_out45 , reg_out46 , reg_out47 , reg_out48 , reg_out49 , reg_out50 , reg_out51 , reg_out52 , reg_out53 , reg_out54 , reg_out55 , reg_out56 , reg_out57 , reg_out58 , reg_out59 , reg_out60 , reg_out61 , reg_out62 , reg_out63 , reg_out64 , reg_out65 , reg_out66 , reg_out67 , reg_out68 , reg_out69 , reg_out70 , reg_out71 , reg_out72 , reg_out73 , reg_out74 , reg_out75 , reg_out76 , reg_out77 , reg_out78 , reg_out79 , reg_out80 , reg_out81 , reg_out82 , reg_out83 , reg_out84 , reg_out85 , reg_out86 , reg_out87 , reg_out88 , reg_out89 , reg_out90 , reg_out91 , reg_out92 , reg_out93 , reg_out94 , reg_out95 , reg_out96 , reg_out97 , reg_out98 , reg_out99 , reg_out100 , reg_out101 , reg_out102 , reg_out103 , reg_out104 , reg_out105 , reg_out106 , reg_out107 , reg_out108 , reg_out109 , reg_out110 , reg_out111 , reg_out112 , reg_out113 , reg_out114 , reg_out115 , reg_out116 , reg_out117 , reg_out118 , reg_out119 , reg_out120 , reg_out121 , reg_out122 , reg_out123 , reg_out124 , reg_out125 , reg_out126 , reg_out127 , reg_out128 , reg_out129 , reg_out130 , reg_out131 , reg_out132 , reg_out133 , reg_out134 , reg_out135 , reg_out136 , reg_out137 , reg_out138 , reg_out139 , reg_out140 , reg_out141 , reg_out142 , reg_out143 , reg_out144 , reg_out145 , reg_out146 , reg_out147 , reg_out148 , reg_out149 , reg_out150 , reg_out151 , reg_out152 , reg_out153 , reg_out154 , reg_out155 , reg_out156 , reg_out157 , reg_out158 , reg_out159 , reg_out160 , reg_out161 , reg_out162 , reg_out163 , reg_out164 , reg_out165 , reg_out166 , reg_out167 , reg_out168 , reg_out169 , reg_out170 , reg_out171 , reg_out172 , reg_out173 , reg_out174 , reg_out175 , reg_out176 , reg_out177 , reg_out178 , reg_out179 , reg_out180 , reg_out181 , reg_out182 , reg_out183 , reg_out184 , reg_out185 , reg_out186 , reg_out187 , reg_out188 , reg_out189 , reg_out190 , reg_out191 , reg_out192 , reg_out193 , reg_out194 , reg_out195 , reg_out196 , reg_out197 , reg_out198 , reg_out199 , reg_out200 , reg_out201 , reg_out202 , reg_out203 , reg_out204 , reg_out205 , reg_out206 , reg_out207 , reg_out208 , reg_out209 , reg_out210 , reg_out211 , reg_out212 , reg_out213 , reg_out214 , reg_out215 , reg_out216 , reg_out217 , reg_out218 , reg_out219 , reg_out220 , reg_out221 , reg_out222 , reg_out223 , reg_out224 , reg_out225 , reg_out226 , reg_out227 , reg_out228 , reg_out229 , reg_out230 , reg_out231 , reg_out232 , reg_out233 , reg_out234 , reg_out235 , reg_out236 , reg_out237 , reg_out238 , reg_out239 , reg_out240 , reg_out241 , reg_out242 , reg_out243 , reg_out244 , reg_out245 , reg_out246 , reg_out247 , reg_out248 , reg_out249 , reg_out250 , reg_out251 , reg_out252 , reg_out253 , reg_out254  ;

always@(posedge clk) begin

    reg_out1  <= in1   ;
    reg_out2  <= in2   ;
    reg_out3  <= in3   ;
    reg_out4  <= in4   ;
    reg_out5  <= in5   ;
    reg_out6  <= in6   ;
    reg_out7  <= in7   ;
    reg_out8  <= in8   ;
    reg_out9  <= in9   ;
    reg_out10  <= in10   ;
    reg_out11  <= in11   ;
    reg_out12  <= in12   ;
    reg_out13  <= in13   ;
    reg_out14  <= in14   ;
    reg_out15  <= in15   ;
    reg_out16  <= in16   ;
    reg_out17  <= in17   ;
    reg_out18  <= in18   ;
    reg_out19  <= in19   ;
    reg_out20  <= in20   ;
    reg_out21  <= in21   ;
    reg_out22  <= in22   ;
    reg_out23  <= in23   ;
    reg_out24  <= in24   ;
    reg_out25  <= in25   ;
    reg_out26  <= in26   ;
    reg_out27  <= in27   ;
    reg_out28  <= in28   ;
    reg_out29  <= in29   ;
    reg_out30  <= in30   ;
    reg_out31  <= in31   ;
    reg_out32  <= in32   ;
    reg_out33  <= in33   ;
    reg_out34  <= in34   ;
    reg_out35  <= in35   ;
    reg_out36  <= in36   ;
    reg_out37  <= in37   ;
    reg_out38  <= in38   ;
    reg_out39  <= in39   ;
    reg_out40  <= in40   ;
    reg_out41  <= in41   ;
    reg_out42  <= in42   ;
    reg_out43  <= in43   ;
    reg_out44  <= in44   ;
    reg_out45  <= in45   ;
    reg_out46  <= in46   ;
    reg_out47  <= in47   ;
    reg_out48  <= in48   ;
    reg_out49  <= in49   ;
    reg_out50  <= in50   ;
    reg_out51  <= in51   ;
    reg_out52  <= in52   ;
    reg_out53  <= in53   ;
    reg_out54  <= in54   ;
    reg_out55  <= in55   ;
    reg_out56  <= in56   ;
    reg_out57  <= in57   ;
    reg_out58  <= in58   ;
    reg_out59  <= in59   ;
    reg_out60  <= in60   ;
    reg_out61  <= in61   ;
    reg_out62  <= in62   ;
    reg_out63  <= in63   ;
    reg_out64  <= in64   ;
    reg_out65  <= in65   ;
    reg_out66  <= in66   ;
    reg_out67  <= in67   ;
    reg_out68  <= in68   ;
    reg_out69  <= in69   ;
    reg_out70  <= in70   ;
    reg_out71  <= in71   ;
    reg_out72  <= in72   ;
    reg_out73  <= in73   ;
    reg_out74  <= in74   ;
    reg_out75  <= in75   ;
    reg_out76  <= in76   ;
    reg_out77  <= in77   ;
    reg_out78  <= in78   ;
    reg_out79  <= in79   ;
    reg_out80  <= in80   ;
    reg_out81  <= in81   ;
    reg_out82  <= in82   ;
    reg_out83  <= in83   ;
    reg_out84  <= in84   ;
    reg_out85  <= in85   ;
    reg_out86  <= in86   ;
    reg_out87  <= in87   ;
    reg_out88  <= in88   ;
    reg_out89  <= in89   ;
    reg_out90  <= in90   ;
    reg_out91  <= in91   ;
    reg_out92  <= in92   ;
    reg_out93  <= in93   ;
    reg_out94  <= in94   ;
    reg_out95  <= in95   ;
    reg_out96  <= in96   ;
    reg_out97  <= in97   ;
    reg_out98  <= in98   ;
    reg_out99  <= in99   ;
    reg_out100  <= in100   ;
    reg_out101  <= in101   ;
    reg_out102  <= in102   ;
    reg_out103  <= in103   ;
    reg_out104  <= in104   ;
    reg_out105  <= in105   ;
    reg_out106  <= in106   ;
    reg_out107  <= in107   ;
    reg_out108  <= in108   ;
    reg_out109  <= in109   ;
    reg_out110  <= in110   ;
    reg_out111  <= in111   ;
    reg_out112  <= in112   ;
    reg_out113  <= in113   ;
    reg_out114  <= in114   ;
    reg_out115  <= in115   ;
    reg_out116  <= in116   ;
    reg_out117  <= in117   ;
    reg_out118  <= in118   ;
    reg_out119  <= in119   ;
    reg_out120  <= in120   ;
    reg_out121  <= in121   ;
    reg_out122  <= in122   ;
    reg_out123  <= in123   ;
    reg_out124  <= in124   ;
    reg_out125  <= in125   ;
    reg_out126  <= in126   ;
    reg_out127  <= in127   ;
    reg_out128  <= in128   ;
    reg_out129  <= in129   ;
    reg_out130  <= in130   ;
    reg_out131  <= in131   ;
    reg_out132  <= in132   ;
    reg_out133  <= in133   ;
    reg_out134  <= in134   ;
    reg_out135  <= in135   ;
    reg_out136  <= in136   ;
    reg_out137  <= in137   ;
    reg_out138  <= in138   ;
    reg_out139  <= in139   ;
    reg_out140  <= in140   ;
    reg_out141  <= in141   ;
    reg_out142  <= in142   ;
    reg_out143  <= in143   ;
    reg_out144  <= in144   ;
    reg_out145  <= in145   ;
    reg_out146  <= in146   ;
    reg_out147  <= in147   ;
    reg_out148  <= in148   ;
    reg_out149  <= in149   ;
    reg_out150  <= in150   ;
    reg_out151  <= in151   ;
    reg_out152  <= in152   ;
    reg_out153  <= in153   ;
    reg_out154  <= in154   ;
    reg_out155  <= in155   ;
    reg_out156  <= in156   ;
    reg_out157  <= in157   ;
    reg_out158  <= in158   ;
    reg_out159  <= in159   ;
    reg_out160  <= in160   ;
    reg_out161  <= in161   ;
    reg_out162  <= in162   ;
    reg_out163  <= in163   ;
    reg_out164  <= in164   ;
    reg_out165  <= in165   ;
    reg_out166  <= in166   ;
    reg_out167  <= in167   ;
    reg_out168  <= in168   ;
    reg_out169  <= in169   ;
    reg_out170  <= in170   ;
    reg_out171  <= in171   ;
    reg_out172  <= in172   ;
    reg_out173  <= in173   ;
    reg_out174  <= in174   ;
    reg_out175  <= in175   ;
    reg_out176  <= in176   ;
    reg_out177  <= in177   ;
    reg_out178  <= in178   ;
    reg_out179  <= in179   ;
    reg_out180  <= in180   ;
    reg_out181  <= in181   ;
    reg_out182  <= in182   ;
    reg_out183  <= in183   ;
    reg_out184  <= in184   ;
    reg_out185  <= in185   ;
    reg_out186  <= in186   ;
    reg_out187  <= in187   ;
    reg_out188  <= in188   ;
    reg_out189  <= in189   ;
    reg_out190  <= in190   ;
    reg_out191  <= in191   ;
    reg_out192  <= in192   ;
    reg_out193  <= in193   ;
    reg_out194  <= in194   ;
    reg_out195  <= in195   ;
    reg_out196  <= in196   ;
    reg_out197  <= in197   ;
    reg_out198  <= in198   ;
    reg_out199  <= in199   ;
    reg_out200  <= in200   ;
    reg_out201  <= in201   ;
    reg_out202  <= in202   ;
    reg_out203  <= in203   ;
    reg_out204  <= in204   ;
    reg_out205  <= in205   ;
    reg_out206  <= in206   ;
    reg_out207  <= in207   ;
    reg_out208  <= in208   ;
    reg_out209  <= in209   ;
    reg_out210  <= in210   ;
    reg_out211  <= in211   ;
    reg_out212  <= in212   ;
    reg_out213  <= in213   ;
    reg_out214  <= in214   ;
    reg_out215  <= in215   ;
    reg_out216  <= in216   ;
    reg_out217  <= in217   ;
    reg_out218  <= in218   ;
    reg_out219  <= in219   ;
    reg_out220  <= in220   ;
    reg_out221  <= in221   ;
    reg_out222  <= in222   ;
    reg_out223  <= in223   ;
    reg_out224  <= in224   ;
    reg_out225  <= in225   ;
    reg_out226  <= in226   ;
    reg_out227  <= in227   ;
    reg_out228  <= in228   ;
    reg_out229  <= in229   ;
    reg_out230  <= in230   ;
    reg_out231  <= in231   ;
    reg_out232  <= in232   ;
    reg_out233  <= in233   ;
    reg_out234  <= in234   ;
    reg_out235  <= in235   ;
    reg_out236  <= in236   ;
    reg_out237  <= in237   ;
    reg_out238  <= in238   ;
    reg_out239  <= in239   ;
    reg_out240  <= in240   ;
    reg_out241  <= in241   ;
    reg_out242  <= in242   ;
    reg_out243  <= in243   ;
    reg_out244  <= in244   ;
    reg_out245  <= in245   ;
    reg_out246  <= in246   ;
    reg_out247  <= in247   ;
    reg_out248  <= in248   ;
    reg_out249  <= in249   ;
    reg_out250  <= in250   ;
    reg_out251  <= in251   ;
    reg_out252  <= in252   ;
    reg_out253  <= in253   ;
    reg_out254  <= in254   ;

end

assign out1 = reg_out1 ;
assign out2 = reg_out2 ;
assign out3 = reg_out3 ;
assign out4 = reg_out4 ;
assign out5 = reg_out5 ;
assign out6 = reg_out6 ;
assign out7 = reg_out7 ;
assign out8 = reg_out8 ;
assign out9 = reg_out9 ;
assign out10 = reg_out10 ;
assign out11 = reg_out11 ;
assign out12 = reg_out12 ;
assign out13 = reg_out13 ;
assign out14 = reg_out14 ;
assign out15 = reg_out15 ;
assign out16 = reg_out16 ;
assign out17 = reg_out17 ;
assign out18 = reg_out18 ;
assign out19 = reg_out19 ;
assign out20 = reg_out20 ;
assign out21 = reg_out21 ;
assign out22 = reg_out22 ;
assign out23 = reg_out23 ;
assign out24 = reg_out24 ;
assign out25 = reg_out25 ;
assign out26 = reg_out26 ;
assign out27 = reg_out27 ;
assign out28 = reg_out28 ;
assign out29 = reg_out29 ;
assign out30 = reg_out30 ;
assign out31 = reg_out31 ;
assign out32 = reg_out32 ;
assign out33 = reg_out33 ;
assign out34 = reg_out34 ;
assign out35 = reg_out35 ;
assign out36 = reg_out36 ;
assign out37 = reg_out37 ;
assign out38 = reg_out38 ;
assign out39 = reg_out39 ;
assign out40 = reg_out40 ;
assign out41 = reg_out41 ;
assign out42 = reg_out42 ;
assign out43 = reg_out43 ;
assign out44 = reg_out44 ;
assign out45 = reg_out45 ;
assign out46 = reg_out46 ;
assign out47 = reg_out47 ;
assign out48 = reg_out48 ;
assign out49 = reg_out49 ;
assign out50 = reg_out50 ;
assign out51 = reg_out51 ;
assign out52 = reg_out52 ;
assign out53 = reg_out53 ;
assign out54 = reg_out54 ;
assign out55 = reg_out55 ;
assign out56 = reg_out56 ;
assign out57 = reg_out57 ;
assign out58 = reg_out58 ;
assign out59 = reg_out59 ;
assign out60 = reg_out60 ;
assign out61 = reg_out61 ;
assign out62 = reg_out62 ;
assign out63 = reg_out63 ;
assign out64 = reg_out64 ;
assign out65 = reg_out65 ;
assign out66 = reg_out66 ;
assign out67 = reg_out67 ;
assign out68 = reg_out68 ;
assign out69 = reg_out69 ;
assign out70 = reg_out70 ;
assign out71 = reg_out71 ;
assign out72 = reg_out72 ;
assign out73 = reg_out73 ;
assign out74 = reg_out74 ;
assign out75 = reg_out75 ;
assign out76 = reg_out76 ;
assign out77 = reg_out77 ;
assign out78 = reg_out78 ;
assign out79 = reg_out79 ;
assign out80 = reg_out80 ;
assign out81 = reg_out81 ;
assign out82 = reg_out82 ;
assign out83 = reg_out83 ;
assign out84 = reg_out84 ;
assign out85 = reg_out85 ;
assign out86 = reg_out86 ;
assign out87 = reg_out87 ;
assign out88 = reg_out88 ;
assign out89 = reg_out89 ;
assign out90 = reg_out90 ;
assign out91 = reg_out91 ;
assign out92 = reg_out92 ;
assign out93 = reg_out93 ;
assign out94 = reg_out94 ;
assign out95 = reg_out95 ;
assign out96 = reg_out96 ;
assign out97 = reg_out97 ;
assign out98 = reg_out98 ;
assign out99 = reg_out99 ;
assign out100 = reg_out100 ;
assign out101 = reg_out101 ;
assign out102 = reg_out102 ;
assign out103 = reg_out103 ;
assign out104 = reg_out104 ;
assign out105 = reg_out105 ;
assign out106 = reg_out106 ;
assign out107 = reg_out107 ;
assign out108 = reg_out108 ;
assign out109 = reg_out109 ;
assign out110 = reg_out110 ;
assign out111 = reg_out111 ;
assign out112 = reg_out112 ;
assign out113 = reg_out113 ;
assign out114 = reg_out114 ;
assign out115 = reg_out115 ;
assign out116 = reg_out116 ;
assign out117 = reg_out117 ;
assign out118 = reg_out118 ;
assign out119 = reg_out119 ;
assign out120 = reg_out120 ;
assign out121 = reg_out121 ;
assign out122 = reg_out122 ;
assign out123 = reg_out123 ;
assign out124 = reg_out124 ;
assign out125 = reg_out125 ;
assign out126 = reg_out126 ;
assign out127 = reg_out127 ;
assign out128 = reg_out128 ;
assign out129 = reg_out129 ;
assign out130 = reg_out130 ;
assign out131 = reg_out131 ;
assign out132 = reg_out132 ;
assign out133 = reg_out133 ;
assign out134 = reg_out134 ;
assign out135 = reg_out135 ;
assign out136 = reg_out136 ;
assign out137 = reg_out137 ;
assign out138 = reg_out138 ;
assign out139 = reg_out139 ;
assign out140 = reg_out140 ;
assign out141 = reg_out141 ;
assign out142 = reg_out142 ;
assign out143 = reg_out143 ;
assign out144 = reg_out144 ;
assign out145 = reg_out145 ;
assign out146 = reg_out146 ;
assign out147 = reg_out147 ;
assign out148 = reg_out148 ;
assign out149 = reg_out149 ;
assign out150 = reg_out150 ;
assign out151 = reg_out151 ;
assign out152 = reg_out152 ;
assign out153 = reg_out153 ;
assign out154 = reg_out154 ;
assign out155 = reg_out155 ;
assign out156 = reg_out156 ;
assign out157 = reg_out157 ;
assign out158 = reg_out158 ;
assign out159 = reg_out159 ;
assign out160 = reg_out160 ;
assign out161 = reg_out161 ;
assign out162 = reg_out162 ;
assign out163 = reg_out163 ;
assign out164 = reg_out164 ;
assign out165 = reg_out165 ;
assign out166 = reg_out166 ;
assign out167 = reg_out167 ;
assign out168 = reg_out168 ;
assign out169 = reg_out169 ;
assign out170 = reg_out170 ;
assign out171 = reg_out171 ;
assign out172 = reg_out172 ;
assign out173 = reg_out173 ;
assign out174 = reg_out174 ;
assign out175 = reg_out175 ;
assign out176 = reg_out176 ;
assign out177 = reg_out177 ;
assign out178 = reg_out178 ;
assign out179 = reg_out179 ;
assign out180 = reg_out180 ;
assign out181 = reg_out181 ;
assign out182 = reg_out182 ;
assign out183 = reg_out183 ;
assign out184 = reg_out184 ;
assign out185 = reg_out185 ;
assign out186 = reg_out186 ;
assign out187 = reg_out187 ;
assign out188 = reg_out188 ;
assign out189 = reg_out189 ;
assign out190 = reg_out190 ;
assign out191 = reg_out191 ;
assign out192 = reg_out192 ;
assign out193 = reg_out193 ;
assign out194 = reg_out194 ;
assign out195 = reg_out195 ;
assign out196 = reg_out196 ;
assign out197 = reg_out197 ;
assign out198 = reg_out198 ;
assign out199 = reg_out199 ;
assign out200 = reg_out200 ;
assign out201 = reg_out201 ;
assign out202 = reg_out202 ;
assign out203 = reg_out203 ;
assign out204 = reg_out204 ;
assign out205 = reg_out205 ;
assign out206 = reg_out206 ;
assign out207 = reg_out207 ;
assign out208 = reg_out208 ;
assign out209 = reg_out209 ;
assign out210 = reg_out210 ;
assign out211 = reg_out211 ;
assign out212 = reg_out212 ;
assign out213 = reg_out213 ;
assign out214 = reg_out214 ;
assign out215 = reg_out215 ;
assign out216 = reg_out216 ;
assign out217 = reg_out217 ;
assign out218 = reg_out218 ;
assign out219 = reg_out219 ;
assign out220 = reg_out220 ;
assign out221 = reg_out221 ;
assign out222 = reg_out222 ;
assign out223 = reg_out223 ;
assign out224 = reg_out224 ;
assign out225 = reg_out225 ;
assign out226 = reg_out226 ;
assign out227 = reg_out227 ;
assign out228 = reg_out228 ;
assign out229 = reg_out229 ;
assign out230 = reg_out230 ;
assign out231 = reg_out231 ;
assign out232 = reg_out232 ;
assign out233 = reg_out233 ;
assign out234 = reg_out234 ;
assign out235 = reg_out235 ;
assign out236 = reg_out236 ;
assign out237 = reg_out237 ;
assign out238 = reg_out238 ;
assign out239 = reg_out239 ;
assign out240 = reg_out240 ;
assign out241 = reg_out241 ;
assign out242 = reg_out242 ;
assign out243 = reg_out243 ;
assign out244 = reg_out244 ;
assign out245 = reg_out245 ;
assign out246 = reg_out246 ;
assign out247 = reg_out247 ;
assign out248 = reg_out248 ;
assign out249 = reg_out249 ;
assign out250 = reg_out250 ;
assign out251 = reg_out251 ;
assign out252 = reg_out252 ;
assign out253 = reg_out253 ;
assign out254 = reg_out254 ;

endmodule