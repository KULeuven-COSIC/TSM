`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper : Time Sharing - A Novel Approach to Low-Latency Masking
// Authors : Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date:    22:18:05 08/23/2023 
// Design Name:    AES S-Box 
// Module Name:    AES_sbox_compute_subscript0 
// Description:    Submodule for AES S-Box. This submodule contains the logic of the first cycle. All crossproducts of the first share.
// 
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module AES_sbox_compute_subscript0( input_share1, rand_bit,  rand_composable_bit,  x0_subscript0_share1_1 , x2_subscript0_share1_1 , x3_subscript0_share1_1 , x4_subscript0_share1_1 , x6_subscript0_share1_1 , x7_subscript0_share1_1 , x1_subscript0_share1_1 , x5_subscript0_share1_1 , x0x1_subscript0_share1_1 , x0x4_subscript0_share1_1 , x0x5_subscript0_share1_1 , x0x6_subscript0_share1_1 , x1x2_subscript0_share1_1 , x1x3_subscript0_share1_1 , x1x4_subscript0_share1_1 , x1x6_subscript0_share1_1 , x2x3_subscript0_share1_1 , x2x4_subscript0_share1_1 , x2x6_subscript0_share1_1 , x2x7_subscript0_share1_1 , x4x6_subscript0_share1_1 , x5x6_subscript0_share1_1 , x5x7_subscript0_share1_1 , x6x7_subscript0_share1_1 , x0x2_subscript0_share1_1 , x0x3_subscript0_share1_1 , x0x7_subscript0_share1_1 , x1x7_subscript0_share1_1 , x3x7_subscript0_share1_1 , x4x5_subscript0_share1_1 , x3x4_subscript0_share1_1 , x4x7_subscript0_share1_1 , x3x6_subscript0_share1_1 , x1x5_subscript0_share1_1 , x2x5_subscript0_share1_1 , x3x5_subscript0_share1_1 , x0x1x4_subscript0_share1_1 , x0x1x6_subscript0_share1_1 , x0x1x7_subscript0_share1_1 , x0x2x4_subscript0_share1_1 , x0x2x5_subscript0_share1_1 , x0x2x6_subscript0_share1_1 , x0x2x7_subscript0_share1_1 , x0x3x4_subscript0_share1_1 , x0x3x5_subscript0_share1_1 , x0x3x6_subscript0_share1_1 , x0x4x6_subscript0_share1_1 , x0x4x7_subscript0_share1_1 , x1x2x3_subscript0_share1_1 , x1x2x4_subscript0_share1_1 , x1x2x6_subscript0_share1_1 , x1x3x4_subscript0_share1_1 , x1x3x7_subscript0_share1_1 , x1x4x6_subscript0_share1_1 , x1x5x6_subscript0_share1_1 , x2x3x5_subscript0_share1_1 , x2x3x7_subscript0_share1_1 , x2x4x7_subscript0_share1_1 , x2x5x6_subscript0_share1_1 , x2x5x7_subscript0_share1_1 , x2x6x7_subscript0_share1_1 , x3x4x7_subscript0_share1_1 , x3x5x7_subscript0_share1_1 , x3x6x7_subscript0_share1_1 , x4x5x6_subscript0_share1_1 , x5x6x7_subscript0_share1_1 , x0x1x3_subscript0_share1_1 , x0x2x3_subscript0_share1_1 , x0x4x5_subscript0_share1_1 , x0x5x7_subscript0_share1_1 , x0x6x7_subscript0_share1_1 , x1x3x5_subscript0_share1_1 , x1x3x6_subscript0_share1_1 , x1x4x7_subscript0_share1_1 , x2x3x4_subscript0_share1_1 , x2x3x6_subscript0_share1_1 , x3x4x6_subscript0_share1_1 , x3x5x6_subscript0_share1_1 , x0x1x5_subscript0_share1_1 , x0x3x7_subscript0_share1_1 , x1x2x5_subscript0_share1_1 , x1x2x7_subscript0_share1_1 , x1x4x5_subscript0_share1_1 , x1x5x7_subscript0_share1_1 , x2x4x5_subscript0_share1_1 , x3x4x5_subscript0_share1_1 , x4x6x7_subscript0_share1_1 , x1x6x7_subscript0_share1_1 , x4x5x7_subscript0_share1_1 , x0x1x2_subscript0_share1_1 , x0x5x6_subscript0_share1_1 , x2x4x6_subscript0_share1_1 , x0x1x2x3_subscript0_share1_1 , x0x1x2x5_subscript0_share1_1 , x0x1x2x6_subscript0_share1_1 , x0x1x2x7_subscript0_share1_1 , x0x1x4x5_subscript0_share1_1 , x0x1x4x7_subscript0_share1_1 , x0x2x3x5_subscript0_share1_1 , x0x2x3x7_subscript0_share1_1 , x0x2x4x5_subscript0_share1_1 , x0x2x4x7_subscript0_share1_1 , x0x2x5x6_subscript0_share1_1 , x0x2x5x7_subscript0_share1_1 , x0x3x4x6_subscript0_share1_1 , x0x3x5x6_subscript0_share1_1 , x0x4x5x6_subscript0_share1_1 , x0x4x5x7_subscript0_share1_1 , x0x4x6x7_subscript0_share1_1 , x1x2x3x5_subscript0_share1_1 , x1x2x3x6_subscript0_share1_1 , x1x2x3x7_subscript0_share1_1 , x1x2x4x6_subscript0_share1_1 , x1x2x4x7_subscript0_share1_1 , x1x2x6x7_subscript0_share1_1 , x1x3x4x6_subscript0_share1_1 , x1x3x6x7_subscript0_share1_1 , x1x4x5x6_subscript0_share1_1 , x1x4x5x7_subscript0_share1_1 , x1x5x6x7_subscript0_share1_1 , x2x3x5x7_subscript0_share1_1 , x2x3x6x7_subscript0_share1_1 , x2x4x5x6_subscript0_share1_1 , x2x4x5x7_subscript0_share1_1 , x3x5x6x7_subscript0_share1_1 , x0x1x3x4_subscript0_share1_1 , x0x1x3x6_subscript0_share1_1 , x0x1x5x6_subscript0_share1_1 , x0x2x3x6_subscript0_share1_1 , x0x3x4x5_subscript0_share1_1 , x1x2x5x6_subscript0_share1_1 , x1x2x5x7_subscript0_share1_1 , x1x3x4x5_subscript0_share1_1 , x1x3x4x7_subscript0_share1_1 , x1x3x5x6_subscript0_share1_1 , x1x3x5x7_subscript0_share1_1 , x1x4x6x7_subscript0_share1_1 , x2x3x4x5_subscript0_share1_1 , x2x3x4x7_subscript0_share1_1 , x2x4x6x7_subscript0_share1_1 , x3x4x5x6_subscript0_share1_1 , x3x4x5x7_subscript0_share1_1 , x3x4x6x7_subscript0_share1_1 , x0x1x3x5_subscript0_share1_1 , x0x1x4x6_subscript0_share1_1 , x0x2x3x4_subscript0_share1_1 , x0x2x4x6_subscript0_share1_1 , x0x3x4x7_subscript0_share1_1 , x0x3x5x7_subscript0_share1_1 , x1x2x3x4_subscript0_share1_1 , x2x3x4x6_subscript0_share1_1 , x2x3x5x6_subscript0_share1_1 , x2x5x6x7_subscript0_share1_1 , x4x5x6x7_subscript0_share1_1 , x0x1x2x4_subscript0_share1_1 , x0x1x6x7_subscript0_share1_1 , x0x2x6x7_subscript0_share1_1 , x0x3x6x7_subscript0_share1_1 , x0x5x6x7_subscript0_share1_1 , x1x2x4x5_subscript0_share1_1 , x0x1x3x7_subscript0_share1_1 , x0x1x5x7_subscript0_share1_1 , x0x1x2x3x4_subscript0_share1_1 , x0x1x2x3x6_subscript0_share1_1 , x0x1x2x3x7_subscript0_share1_1 , x0x1x2x4x5_subscript0_share1_1 , x0x1x2x4x7_subscript0_share1_1 , x0x1x2x5x7_subscript0_share1_1 , x0x1x2x6x7_subscript0_share1_1 , x0x1x3x4x6_subscript0_share1_1 , x0x1x3x5x6_subscript0_share1_1 , x0x1x3x5x7_subscript0_share1_1 , x0x1x3x6x7_subscript0_share1_1 , x0x1x4x5x6_subscript0_share1_1 , x0x1x5x6x7_subscript0_share1_1 , x0x2x3x4x5_subscript0_share1_1 , x0x2x3x4x6_subscript0_share1_1 , x0x2x4x5x7_subscript0_share1_1 , x0x2x4x6x7_subscript0_share1_1 , x0x3x4x5x6_subscript0_share1_1 , x0x3x4x5x7_subscript0_share1_1 , x0x3x4x6x7_subscript0_share1_1 , x0x3x5x6x7_subscript0_share1_1 , x1x2x3x5x6_subscript0_share1_1 , x1x2x3x5x7_subscript0_share1_1 , x1x2x4x5x6_subscript0_share1_1 , x1x2x4x6x7_subscript0_share1_1 , x1x2x5x6x7_subscript0_share1_1 , x1x3x4x5x7_subscript0_share1_1 , x2x3x4x5x6_subscript0_share1_1 , x2x3x4x5x7_subscript0_share1_1 , x2x4x5x6x7_subscript0_share1_1 , x0x1x2x4x6_subscript0_share1_1 , x0x1x3x4x7_subscript0_share1_1 , x0x2x3x4x7_subscript0_share1_1 , x0x2x3x5x7_subscript0_share1_1 , x0x2x3x6x7_subscript0_share1_1 , x0x2x4x5x6_subscript0_share1_1 , x0x2x5x6x7_subscript0_share1_1 , x0x4x5x6x7_subscript0_share1_1 , x1x2x3x4x6_subscript0_share1_1 , x1x3x4x5x6_subscript0_share1_1 , x2x3x4x6x7_subscript0_share1_1 , x0x1x2x3x5_subscript0_share1_1 , x0x1x4x6x7_subscript0_share1_1 , x1x2x3x4x5_subscript0_share1_1 , x1x2x3x6x7_subscript0_share1_1 , x1x2x4x5x7_subscript0_share1_1 , x1x3x4x6x7_subscript0_share1_1 , x1x3x5x6x7_subscript0_share1_1 , x1x4x5x6x7_subscript0_share1_1 , x2x3x5x6x7_subscript0_share1_1 , x3x4x5x6x7_subscript0_share1_1 , x0x1x2x5x6_subscript0_share1_1 , x0x1x3x4x5_subscript0_share1_1 , x0x1x4x5x7_subscript0_share1_1 , x0x2x3x5x6_subscript0_share1_1 , x1x2x3x4x7_subscript0_share1_1 , x0x1x2x3x4x6_subscript0_share1_1 , x0x1x2x3x4x7_subscript0_share1_1 , x0x1x2x3x5x7_subscript0_share1_1 , x0x1x2x3x6x7_subscript0_share1_1 , x0x1x2x4x5x7_subscript0_share1_1 , x0x1x2x5x6x7_subscript0_share1_1 , x0x1x3x4x6x7_subscript0_share1_1 , x0x1x4x5x6x7_subscript0_share1_1 , x0x2x3x4x5x6_subscript0_share1_1 , x0x2x3x4x5x7_subscript0_share1_1 , x0x2x3x5x6x7_subscript0_share1_1 , x1x2x3x4x6x7_subscript0_share1_1 , x1x2x4x5x6x7_subscript0_share1_1 , x1x3x4x5x6x7_subscript0_share1_1 , x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x5x6_subscript0_share1_1 , x0x1x2x4x6x7_subscript0_share1_1 , x0x1x3x4x5x6_subscript0_share1_1 , x0x2x3x4x6x7_subscript0_share1_1 , x1x2x3x4x5x6_subscript0_share1_1 , x1x2x3x5x6x7_subscript0_share1_1 , x0x1x2x3x4x5_subscript0_share1_1 , x0x1x2x4x5x6_subscript0_share1_1 , x0x1x3x4x5x7_subscript0_share1_1 , x0x1x3x5x6x7_subscript0_share1_1 , x0x2x4x5x6x7_subscript0_share1_1 , x1x2x3x4x5x7_subscript0_share1_1 , x0x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x4x6x7_subscript0_share1_1 , x0x1x2x4x5x6x7_subscript0_share1_1 , x0x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x5x6x7_subscript0_share1_1 , x0x1x3x4x5x6x7_subscript0_share1_1 , x1x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x4x5x6_subscript0_share1_1 , x0x1x2x3x4x5x7_subscript0_share1_1 , x0_subscript0_share2_1 , x2_subscript0_share2_1 , x3_subscript0_share2_1 , x4_subscript0_share2_1 , x6_subscript0_share2_1 , x7_subscript0_share2_1 , x1_subscript0_share2_1 , x5_subscript0_share2_1 , x0x1_subscript0_share2_1 , x0x4_subscript0_share2_1 , x0x5_subscript0_share2_1 , x0x6_subscript0_share2_1 , x1x2_subscript0_share2_1 , x1x3_subscript0_share2_1 , x1x4_subscript0_share2_1 , x1x6_subscript0_share2_1 , x2x3_subscript0_share2_1 , x2x4_subscript0_share2_1 , x2x6_subscript0_share2_1 , x2x7_subscript0_share2_1 , x4x6_subscript0_share2_1 , x5x6_subscript0_share2_1 , x5x7_subscript0_share2_1 , x6x7_subscript0_share2_1 , x0x2_subscript0_share2_1 , x0x3_subscript0_share2_1 , x0x7_subscript0_share2_1 , x1x7_subscript0_share2_1 , x3x7_subscript0_share2_1 , x4x5_subscript0_share2_1 , x3x4_subscript0_share2_1 , x4x7_subscript0_share2_1 , x3x6_subscript0_share2_1 , x1x5_subscript0_share2_1 , x2x5_subscript0_share2_1 , x3x5_subscript0_share2_1 , x0x1x4_subscript0_share2_1 , x0x1x6_subscript0_share2_1 , x0x1x7_subscript0_share2_1 , x0x2x4_subscript0_share2_1 , x0x2x5_subscript0_share2_1 , x0x2x6_subscript0_share2_1 , x0x2x7_subscript0_share2_1 , x0x3x4_subscript0_share2_1 , x0x3x5_subscript0_share2_1 , x0x3x6_subscript0_share2_1 , x0x4x6_subscript0_share2_1 , x0x4x7_subscript0_share2_1 , x1x2x3_subscript0_share2_1 , x1x2x4_subscript0_share2_1 , x1x2x6_subscript0_share2_1 , x1x3x4_subscript0_share2_1 , x1x3x7_subscript0_share2_1 , x1x4x6_subscript0_share2_1 , x1x5x6_subscript0_share2_1 , x2x3x5_subscript0_share2_1 , x2x3x7_subscript0_share2_1 , x2x4x7_subscript0_share2_1 , x2x5x6_subscript0_share2_1 , x2x5x7_subscript0_share2_1 , x2x6x7_subscript0_share2_1 , x3x4x7_subscript0_share2_1 , x3x5x7_subscript0_share2_1 , x3x6x7_subscript0_share2_1 , x4x5x6_subscript0_share2_1 , x5x6x7_subscript0_share2_1 , x0x1x3_subscript0_share2_1 , x0x2x3_subscript0_share2_1 , x0x4x5_subscript0_share2_1 , x0x5x7_subscript0_share2_1 , x0x6x7_subscript0_share2_1 , x1x3x5_subscript0_share2_1 , x1x3x6_subscript0_share2_1 , x1x4x7_subscript0_share2_1 , x2x3x4_subscript0_share2_1 , x2x3x6_subscript0_share2_1 , x3x4x6_subscript0_share2_1 , x3x5x6_subscript0_share2_1 , x0x1x5_subscript0_share2_1 , x0x3x7_subscript0_share2_1 , x1x2x5_subscript0_share2_1 , x1x2x7_subscript0_share2_1 , x1x4x5_subscript0_share2_1 , x1x5x7_subscript0_share2_1 , x2x4x5_subscript0_share2_1 , x3x4x5_subscript0_share2_1 , x4x6x7_subscript0_share2_1 , x1x6x7_subscript0_share2_1 , x4x5x7_subscript0_share2_1 , x0x1x2_subscript0_share2_1 , x0x5x6_subscript0_share2_1 , x2x4x6_subscript0_share2_1 , x0x1x2x3_subscript0_share2_1 , x0x1x2x5_subscript0_share2_1 , x0x1x2x6_subscript0_share2_1 , x0x1x2x7_subscript0_share2_1 , x0x1x4x5_subscript0_share2_1 , x0x1x4x7_subscript0_share2_1 , x0x2x3x5_subscript0_share2_1 , x0x2x3x7_subscript0_share2_1 , x0x2x4x5_subscript0_share2_1 , x0x2x4x7_subscript0_share2_1 , x0x2x5x6_subscript0_share2_1 , x0x2x5x7_subscript0_share2_1 , x0x3x4x6_subscript0_share2_1 , x0x3x5x6_subscript0_share2_1 , x0x4x5x6_subscript0_share2_1 , x0x4x5x7_subscript0_share2_1 , x0x4x6x7_subscript0_share2_1 , x1x2x3x5_subscript0_share2_1 , x1x2x3x6_subscript0_share2_1 , x1x2x3x7_subscript0_share2_1 , x1x2x4x6_subscript0_share2_1 , x1x2x4x7_subscript0_share2_1 , x1x2x6x7_subscript0_share2_1 , x1x3x4x6_subscript0_share2_1 , x1x3x6x7_subscript0_share2_1 , x1x4x5x6_subscript0_share2_1 , x1x4x5x7_subscript0_share2_1 , x1x5x6x7_subscript0_share2_1 , x2x3x5x7_subscript0_share2_1 , x2x3x6x7_subscript0_share2_1 , x2x4x5x6_subscript0_share2_1 , x2x4x5x7_subscript0_share2_1 , x3x5x6x7_subscript0_share2_1 , x0x1x3x4_subscript0_share2_1 , x0x1x3x6_subscript0_share2_1 , x0x1x5x6_subscript0_share2_1 , x0x2x3x6_subscript0_share2_1 , x0x3x4x5_subscript0_share2_1 , x1x2x5x6_subscript0_share2_1 , x1x2x5x7_subscript0_share2_1 , x1x3x4x5_subscript0_share2_1 , x1x3x4x7_subscript0_share2_1 , x1x3x5x6_subscript0_share2_1 , x1x3x5x7_subscript0_share2_1 , x1x4x6x7_subscript0_share2_1 , x2x3x4x5_subscript0_share2_1 , x2x3x4x7_subscript0_share2_1 , x2x4x6x7_subscript0_share2_1 , x3x4x5x6_subscript0_share2_1 , x3x4x5x7_subscript0_share2_1 , x3x4x6x7_subscript0_share2_1 , x0x1x3x5_subscript0_share2_1 , x0x1x4x6_subscript0_share2_1 , x0x2x3x4_subscript0_share2_1 , x0x2x4x6_subscript0_share2_1 , x0x3x4x7_subscript0_share2_1 , x0x3x5x7_subscript0_share2_1 , x1x2x3x4_subscript0_share2_1 , x2x3x4x6_subscript0_share2_1 , x2x3x5x6_subscript0_share2_1 , x2x5x6x7_subscript0_share2_1 , x4x5x6x7_subscript0_share2_1 , x0x1x2x4_subscript0_share2_1 , x0x1x6x7_subscript0_share2_1 , x0x2x6x7_subscript0_share2_1 , x0x3x6x7_subscript0_share2_1 , x0x5x6x7_subscript0_share2_1 , x1x2x4x5_subscript0_share2_1 , x0x1x3x7_subscript0_share2_1 , x0x1x5x7_subscript0_share2_1 , x0x1x2x3x4_subscript0_share2_1 , x0x1x2x3x6_subscript0_share2_1 , x0x1x2x3x7_subscript0_share2_1 , x0x1x2x4x5_subscript0_share2_1 , x0x1x2x4x7_subscript0_share2_1 , x0x1x2x5x7_subscript0_share2_1 , x0x1x2x6x7_subscript0_share2_1 , x0x1x3x4x6_subscript0_share2_1 , x0x1x3x5x6_subscript0_share2_1 , x0x1x3x5x7_subscript0_share2_1 , x0x1x3x6x7_subscript0_share2_1 , x0x1x4x5x6_subscript0_share2_1 , x0x1x5x6x7_subscript0_share2_1 , x0x2x3x4x5_subscript0_share2_1 , x0x2x3x4x6_subscript0_share2_1 , x0x2x4x5x7_subscript0_share2_1 , x0x2x4x6x7_subscript0_share2_1 , x0x3x4x5x6_subscript0_share2_1 , x0x3x4x5x7_subscript0_share2_1 , x0x3x4x6x7_subscript0_share2_1 , x0x3x5x6x7_subscript0_share2_1 , x1x2x3x5x6_subscript0_share2_1 , x1x2x3x5x7_subscript0_share2_1 , x1x2x4x5x6_subscript0_share2_1 , x1x2x4x6x7_subscript0_share2_1 , x1x2x5x6x7_subscript0_share2_1 , x1x3x4x5x7_subscript0_share2_1 , x2x3x4x5x6_subscript0_share2_1 , x2x3x4x5x7_subscript0_share2_1 , x2x4x5x6x7_subscript0_share2_1 , x0x1x2x4x6_subscript0_share2_1 , x0x1x3x4x7_subscript0_share2_1 , x0x2x3x4x7_subscript0_share2_1 , x0x2x3x5x7_subscript0_share2_1 , x0x2x3x6x7_subscript0_share2_1 , x0x2x4x5x6_subscript0_share2_1 , x0x2x5x6x7_subscript0_share2_1 , x0x4x5x6x7_subscript0_share2_1 , x1x2x3x4x6_subscript0_share2_1 , x1x3x4x5x6_subscript0_share2_1 , x2x3x4x6x7_subscript0_share2_1 , x0x1x2x3x5_subscript0_share2_1 , x0x1x4x6x7_subscript0_share2_1 , x1x2x3x4x5_subscript0_share2_1 , x1x2x3x6x7_subscript0_share2_1 , x1x2x4x5x7_subscript0_share2_1 , x1x3x4x6x7_subscript0_share2_1 , x1x3x5x6x7_subscript0_share2_1 , x1x4x5x6x7_subscript0_share2_1 , x2x3x5x6x7_subscript0_share2_1 , x3x4x5x6x7_subscript0_share2_1 , x0x1x2x5x6_subscript0_share2_1 , x0x1x3x4x5_subscript0_share2_1 , x0x1x4x5x7_subscript0_share2_1 , x0x2x3x5x6_subscript0_share2_1 , x1x2x3x4x7_subscript0_share2_1 , x0x1x2x3x4x6_subscript0_share2_1 , x0x1x2x3x4x7_subscript0_share2_1 , x0x1x2x3x5x7_subscript0_share2_1 , x0x1x2x3x6x7_subscript0_share2_1 , x0x1x2x4x5x7_subscript0_share2_1 , x0x1x2x5x6x7_subscript0_share2_1 , x0x1x3x4x6x7_subscript0_share2_1 , x0x1x4x5x6x7_subscript0_share2_1 , x0x2x3x4x5x6_subscript0_share2_1 , x0x2x3x4x5x7_subscript0_share2_1 , x0x2x3x5x6x7_subscript0_share2_1 , x1x2x3x4x6x7_subscript0_share2_1 , x1x2x4x5x6x7_subscript0_share2_1 , x1x3x4x5x6x7_subscript0_share2_1 , x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x5x6_subscript0_share2_1 , x0x1x2x4x6x7_subscript0_share2_1 , x0x1x3x4x5x6_subscript0_share2_1 , x0x2x3x4x6x7_subscript0_share2_1 , x1x2x3x4x5x6_subscript0_share2_1 , x1x2x3x5x6x7_subscript0_share2_1 , x0x1x2x3x4x5_subscript0_share2_1 , x0x1x2x4x5x6_subscript0_share2_1 , x0x1x3x4x5x7_subscript0_share2_1 , x0x1x3x5x6x7_subscript0_share2_1 , x0x2x4x5x6x7_subscript0_share2_1 , x1x2x3x4x5x7_subscript0_share2_1 , x0x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x4x6x7_subscript0_share2_1 , x0x1x2x4x5x6x7_subscript0_share2_1 , x0x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x5x6x7_subscript0_share2_1 , x0x1x3x4x5x6x7_subscript0_share2_1 , x1x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x4x5x6_subscript0_share2_1 , x0x1x2x3x4x5x7_subscript0_share2_1 );

input [7:0] input_share1 ;
input [254:1] rand_bit ;
input [7:0] rand_composable_bit ;

output x0_subscript0_share1_1 , x2_subscript0_share1_1 , x3_subscript0_share1_1 , x4_subscript0_share1_1 , x6_subscript0_share1_1 , x7_subscript0_share1_1 , x1_subscript0_share1_1 , x5_subscript0_share1_1 , x0x1_subscript0_share1_1 , x0x4_subscript0_share1_1 , x0x5_subscript0_share1_1 , x0x6_subscript0_share1_1 , x1x2_subscript0_share1_1 , x1x3_subscript0_share1_1 , x1x4_subscript0_share1_1 , x1x6_subscript0_share1_1 , x2x3_subscript0_share1_1 , x2x4_subscript0_share1_1 , x2x6_subscript0_share1_1 , x2x7_subscript0_share1_1 , x4x6_subscript0_share1_1 , x5x6_subscript0_share1_1 , x5x7_subscript0_share1_1 , x6x7_subscript0_share1_1 , x0x2_subscript0_share1_1 , x0x3_subscript0_share1_1 , x0x7_subscript0_share1_1 , x1x7_subscript0_share1_1 , x3x7_subscript0_share1_1 , x4x5_subscript0_share1_1 , x3x4_subscript0_share1_1 , x4x7_subscript0_share1_1 , x3x6_subscript0_share1_1 , x1x5_subscript0_share1_1 , x2x5_subscript0_share1_1 , x3x5_subscript0_share1_1 , x0x1x4_subscript0_share1_1 , x0x1x6_subscript0_share1_1 , x0x1x7_subscript0_share1_1 , x0x2x4_subscript0_share1_1 , x0x2x5_subscript0_share1_1 , x0x2x6_subscript0_share1_1 , x0x2x7_subscript0_share1_1 , x0x3x4_subscript0_share1_1 , x0x3x5_subscript0_share1_1 , x0x3x6_subscript0_share1_1 , x0x4x6_subscript0_share1_1 , x0x4x7_subscript0_share1_1 , x1x2x3_subscript0_share1_1 , x1x2x4_subscript0_share1_1 , x1x2x6_subscript0_share1_1 , x1x3x4_subscript0_share1_1 , x1x3x7_subscript0_share1_1 , x1x4x6_subscript0_share1_1 , x1x5x6_subscript0_share1_1 , x2x3x5_subscript0_share1_1 , x2x3x7_subscript0_share1_1 , x2x4x7_subscript0_share1_1 , x2x5x6_subscript0_share1_1 , x2x5x7_subscript0_share1_1 , x2x6x7_subscript0_share1_1 , x3x4x7_subscript0_share1_1 , x3x5x7_subscript0_share1_1 , x3x6x7_subscript0_share1_1 , x4x5x6_subscript0_share1_1 , x5x6x7_subscript0_share1_1 , x0x1x3_subscript0_share1_1 , x0x2x3_subscript0_share1_1 , x0x4x5_subscript0_share1_1 , x0x5x7_subscript0_share1_1 , x0x6x7_subscript0_share1_1 , x1x3x5_subscript0_share1_1 , x1x3x6_subscript0_share1_1 , x1x4x7_subscript0_share1_1 , x2x3x4_subscript0_share1_1 , x2x3x6_subscript0_share1_1 , x3x4x6_subscript0_share1_1 , x3x5x6_subscript0_share1_1 , x0x1x5_subscript0_share1_1 , x0x3x7_subscript0_share1_1 , x1x2x5_subscript0_share1_1 , x1x2x7_subscript0_share1_1 , x1x4x5_subscript0_share1_1 , x1x5x7_subscript0_share1_1 , x2x4x5_subscript0_share1_1 , x3x4x5_subscript0_share1_1 , x4x6x7_subscript0_share1_1 , x1x6x7_subscript0_share1_1 , x4x5x7_subscript0_share1_1 , x0x1x2_subscript0_share1_1 , x0x5x6_subscript0_share1_1 , x2x4x6_subscript0_share1_1 , x0x1x2x3_subscript0_share1_1 , x0x1x2x5_subscript0_share1_1 , x0x1x2x6_subscript0_share1_1 , x0x1x2x7_subscript0_share1_1 , x0x1x4x5_subscript0_share1_1 , x0x1x4x7_subscript0_share1_1 , x0x2x3x5_subscript0_share1_1 , x0x2x3x7_subscript0_share1_1 , x0x2x4x5_subscript0_share1_1 , x0x2x4x7_subscript0_share1_1 , x0x2x5x6_subscript0_share1_1 , x0x2x5x7_subscript0_share1_1 , x0x3x4x6_subscript0_share1_1 , x0x3x5x6_subscript0_share1_1 , x0x4x5x6_subscript0_share1_1 , x0x4x5x7_subscript0_share1_1 , x0x4x6x7_subscript0_share1_1 , x1x2x3x5_subscript0_share1_1 , x1x2x3x6_subscript0_share1_1 , x1x2x3x7_subscript0_share1_1 , x1x2x4x6_subscript0_share1_1 , x1x2x4x7_subscript0_share1_1 , x1x2x6x7_subscript0_share1_1 , x1x3x4x6_subscript0_share1_1 , x1x3x6x7_subscript0_share1_1 , x1x4x5x6_subscript0_share1_1 , x1x4x5x7_subscript0_share1_1 , x1x5x6x7_subscript0_share1_1 , x2x3x5x7_subscript0_share1_1 , x2x3x6x7_subscript0_share1_1 , x2x4x5x6_subscript0_share1_1 , x2x4x5x7_subscript0_share1_1 , x3x5x6x7_subscript0_share1_1 , x0x1x3x4_subscript0_share1_1 , x0x1x3x6_subscript0_share1_1 , x0x1x5x6_subscript0_share1_1 , x0x2x3x6_subscript0_share1_1 , x0x3x4x5_subscript0_share1_1 , x1x2x5x6_subscript0_share1_1 , x1x2x5x7_subscript0_share1_1 , x1x3x4x5_subscript0_share1_1 , x1x3x4x7_subscript0_share1_1 , x1x3x5x6_subscript0_share1_1 , x1x3x5x7_subscript0_share1_1 , x1x4x6x7_subscript0_share1_1 , x2x3x4x5_subscript0_share1_1 , x2x3x4x7_subscript0_share1_1 , x2x4x6x7_subscript0_share1_1 , x3x4x5x6_subscript0_share1_1 , x3x4x5x7_subscript0_share1_1 , x3x4x6x7_subscript0_share1_1 , x0x1x3x5_subscript0_share1_1 , x0x1x4x6_subscript0_share1_1 , x0x2x3x4_subscript0_share1_1 , x0x2x4x6_subscript0_share1_1 , x0x3x4x7_subscript0_share1_1 , x0x3x5x7_subscript0_share1_1 , x1x2x3x4_subscript0_share1_1 , x2x3x4x6_subscript0_share1_1 , x2x3x5x6_subscript0_share1_1 , x2x5x6x7_subscript0_share1_1 , x4x5x6x7_subscript0_share1_1 , x0x1x2x4_subscript0_share1_1 , x0x1x6x7_subscript0_share1_1 , x0x2x6x7_subscript0_share1_1 , x0x3x6x7_subscript0_share1_1 , x0x5x6x7_subscript0_share1_1 , x1x2x4x5_subscript0_share1_1 , x0x1x3x7_subscript0_share1_1 , x0x1x5x7_subscript0_share1_1 , x0x1x2x3x4_subscript0_share1_1 , x0x1x2x3x6_subscript0_share1_1 , x0x1x2x3x7_subscript0_share1_1 , x0x1x2x4x5_subscript0_share1_1 , x0x1x2x4x7_subscript0_share1_1 , x0x1x2x5x7_subscript0_share1_1 , x0x1x2x6x7_subscript0_share1_1 , x0x1x3x4x6_subscript0_share1_1 , x0x1x3x5x6_subscript0_share1_1 , x0x1x3x5x7_subscript0_share1_1 , x0x1x3x6x7_subscript0_share1_1 , x0x1x4x5x6_subscript0_share1_1 , x0x1x5x6x7_subscript0_share1_1 , x0x2x3x4x5_subscript0_share1_1 , x0x2x3x4x6_subscript0_share1_1 , x0x2x4x5x7_subscript0_share1_1 , x0x2x4x6x7_subscript0_share1_1 , x0x3x4x5x6_subscript0_share1_1 , x0x3x4x5x7_subscript0_share1_1 , x0x3x4x6x7_subscript0_share1_1 , x0x3x5x6x7_subscript0_share1_1 , x1x2x3x5x6_subscript0_share1_1 , x1x2x3x5x7_subscript0_share1_1 , x1x2x4x5x6_subscript0_share1_1 , x1x2x4x6x7_subscript0_share1_1 , x1x2x5x6x7_subscript0_share1_1 , x1x3x4x5x7_subscript0_share1_1 , x2x3x4x5x6_subscript0_share1_1 , x2x3x4x5x7_subscript0_share1_1 , x2x4x5x6x7_subscript0_share1_1 , x0x1x2x4x6_subscript0_share1_1 , x0x1x3x4x7_subscript0_share1_1 , x0x2x3x4x7_subscript0_share1_1 , x0x2x3x5x7_subscript0_share1_1 , x0x2x3x6x7_subscript0_share1_1 , x0x2x4x5x6_subscript0_share1_1 , x0x2x5x6x7_subscript0_share1_1 , x0x4x5x6x7_subscript0_share1_1 , x1x2x3x4x6_subscript0_share1_1 , x1x3x4x5x6_subscript0_share1_1 , x2x3x4x6x7_subscript0_share1_1 , x0x1x2x3x5_subscript0_share1_1 , x0x1x4x6x7_subscript0_share1_1 , x1x2x3x4x5_subscript0_share1_1 , x1x2x3x6x7_subscript0_share1_1 , x1x2x4x5x7_subscript0_share1_1 , x1x3x4x6x7_subscript0_share1_1 , x1x3x5x6x7_subscript0_share1_1 , x1x4x5x6x7_subscript0_share1_1 , x2x3x5x6x7_subscript0_share1_1 , x3x4x5x6x7_subscript0_share1_1 , x0x1x2x5x6_subscript0_share1_1 , x0x1x3x4x5_subscript0_share1_1 , x0x1x4x5x7_subscript0_share1_1 , x0x2x3x5x6_subscript0_share1_1 , x1x2x3x4x7_subscript0_share1_1 , x0x1x2x3x4x6_subscript0_share1_1 , x0x1x2x3x4x7_subscript0_share1_1 , x0x1x2x3x5x7_subscript0_share1_1 , x0x1x2x3x6x7_subscript0_share1_1 , x0x1x2x4x5x7_subscript0_share1_1 , x0x1x2x5x6x7_subscript0_share1_1 , x0x1x3x4x6x7_subscript0_share1_1 , x0x1x4x5x6x7_subscript0_share1_1 , x0x2x3x4x5x6_subscript0_share1_1 , x0x2x3x4x5x7_subscript0_share1_1 , x0x2x3x5x6x7_subscript0_share1_1 , x1x2x3x4x6x7_subscript0_share1_1 , x1x2x4x5x6x7_subscript0_share1_1 , x1x3x4x5x6x7_subscript0_share1_1 , x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x5x6_subscript0_share1_1 , x0x1x2x4x6x7_subscript0_share1_1 , x0x1x3x4x5x6_subscript0_share1_1 , x0x2x3x4x6x7_subscript0_share1_1 , x1x2x3x4x5x6_subscript0_share1_1 , x1x2x3x5x6x7_subscript0_share1_1 , x0x1x2x3x4x5_subscript0_share1_1 , x0x1x2x4x5x6_subscript0_share1_1 , x0x1x3x4x5x7_subscript0_share1_1 , x0x1x3x5x6x7_subscript0_share1_1 , x0x2x4x5x6x7_subscript0_share1_1 , x1x2x3x4x5x7_subscript0_share1_1 , x0x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x4x6x7_subscript0_share1_1 , x0x1x2x4x5x6x7_subscript0_share1_1 , x0x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x5x6x7_subscript0_share1_1 , x0x1x3x4x5x6x7_subscript0_share1_1 , x1x2x3x4x5x6x7_subscript0_share1_1 , x0x1x2x3x4x5x6_subscript0_share1_1 , x0x1x2x3x4x5x7_subscript0_share1_1 , x0_subscript0_share2_1 , x2_subscript0_share2_1 , x3_subscript0_share2_1 , x4_subscript0_share2_1 , x6_subscript0_share2_1 , x7_subscript0_share2_1 , x1_subscript0_share2_1 , x5_subscript0_share2_1 , x0x1_subscript0_share2_1 , x0x4_subscript0_share2_1 , x0x5_subscript0_share2_1 , x0x6_subscript0_share2_1 , x1x2_subscript0_share2_1 , x1x3_subscript0_share2_1 , x1x4_subscript0_share2_1 , x1x6_subscript0_share2_1 , x2x3_subscript0_share2_1 , x2x4_subscript0_share2_1 , x2x6_subscript0_share2_1 , x2x7_subscript0_share2_1 , x4x6_subscript0_share2_1 , x5x6_subscript0_share2_1 , x5x7_subscript0_share2_1 , x6x7_subscript0_share2_1 , x0x2_subscript0_share2_1 , x0x3_subscript0_share2_1 , x0x7_subscript0_share2_1 , x1x7_subscript0_share2_1 , x3x7_subscript0_share2_1 , x4x5_subscript0_share2_1 , x3x4_subscript0_share2_1 , x4x7_subscript0_share2_1 , x3x6_subscript0_share2_1 , x1x5_subscript0_share2_1 , x2x5_subscript0_share2_1 , x3x5_subscript0_share2_1 , x0x1x4_subscript0_share2_1 , x0x1x6_subscript0_share2_1 , x0x1x7_subscript0_share2_1 , x0x2x4_subscript0_share2_1 , x0x2x5_subscript0_share2_1 , x0x2x6_subscript0_share2_1 , x0x2x7_subscript0_share2_1 , x0x3x4_subscript0_share2_1 , x0x3x5_subscript0_share2_1 , x0x3x6_subscript0_share2_1 , x0x4x6_subscript0_share2_1 , x0x4x7_subscript0_share2_1 , x1x2x3_subscript0_share2_1 , x1x2x4_subscript0_share2_1 , x1x2x6_subscript0_share2_1 , x1x3x4_subscript0_share2_1 , x1x3x7_subscript0_share2_1 , x1x4x6_subscript0_share2_1 , x1x5x6_subscript0_share2_1 , x2x3x5_subscript0_share2_1 , x2x3x7_subscript0_share2_1 , x2x4x7_subscript0_share2_1 , x2x5x6_subscript0_share2_1 , x2x5x7_subscript0_share2_1 , x2x6x7_subscript0_share2_1 , x3x4x7_subscript0_share2_1 , x3x5x7_subscript0_share2_1 , x3x6x7_subscript0_share2_1 , x4x5x6_subscript0_share2_1 , x5x6x7_subscript0_share2_1 , x0x1x3_subscript0_share2_1 , x0x2x3_subscript0_share2_1 , x0x4x5_subscript0_share2_1 , x0x5x7_subscript0_share2_1 , x0x6x7_subscript0_share2_1 , x1x3x5_subscript0_share2_1 , x1x3x6_subscript0_share2_1 , x1x4x7_subscript0_share2_1 , x2x3x4_subscript0_share2_1 , x2x3x6_subscript0_share2_1 , x3x4x6_subscript0_share2_1 , x3x5x6_subscript0_share2_1 , x0x1x5_subscript0_share2_1 , x0x3x7_subscript0_share2_1 , x1x2x5_subscript0_share2_1 , x1x2x7_subscript0_share2_1 , x1x4x5_subscript0_share2_1 , x1x5x7_subscript0_share2_1 , x2x4x5_subscript0_share2_1 , x3x4x5_subscript0_share2_1 , x4x6x7_subscript0_share2_1 , x1x6x7_subscript0_share2_1 , x4x5x7_subscript0_share2_1 , x0x1x2_subscript0_share2_1 , x0x5x6_subscript0_share2_1 , x2x4x6_subscript0_share2_1 , x0x1x2x3_subscript0_share2_1 , x0x1x2x5_subscript0_share2_1 , x0x1x2x6_subscript0_share2_1 , x0x1x2x7_subscript0_share2_1 , x0x1x4x5_subscript0_share2_1 , x0x1x4x7_subscript0_share2_1 , x0x2x3x5_subscript0_share2_1 , x0x2x3x7_subscript0_share2_1 , x0x2x4x5_subscript0_share2_1 , x0x2x4x7_subscript0_share2_1 , x0x2x5x6_subscript0_share2_1 , x0x2x5x7_subscript0_share2_1 , x0x3x4x6_subscript0_share2_1 , x0x3x5x6_subscript0_share2_1 , x0x4x5x6_subscript0_share2_1 , x0x4x5x7_subscript0_share2_1 , x0x4x6x7_subscript0_share2_1 , x1x2x3x5_subscript0_share2_1 , x1x2x3x6_subscript0_share2_1 , x1x2x3x7_subscript0_share2_1 , x1x2x4x6_subscript0_share2_1 , x1x2x4x7_subscript0_share2_1 , x1x2x6x7_subscript0_share2_1 , x1x3x4x6_subscript0_share2_1 , x1x3x6x7_subscript0_share2_1 , x1x4x5x6_subscript0_share2_1 , x1x4x5x7_subscript0_share2_1 , x1x5x6x7_subscript0_share2_1 , x2x3x5x7_subscript0_share2_1 , x2x3x6x7_subscript0_share2_1 , x2x4x5x6_subscript0_share2_1 , x2x4x5x7_subscript0_share2_1 , x3x5x6x7_subscript0_share2_1 , x0x1x3x4_subscript0_share2_1 , x0x1x3x6_subscript0_share2_1 , x0x1x5x6_subscript0_share2_1 , x0x2x3x6_subscript0_share2_1 , x0x3x4x5_subscript0_share2_1 , x1x2x5x6_subscript0_share2_1 , x1x2x5x7_subscript0_share2_1 , x1x3x4x5_subscript0_share2_1 , x1x3x4x7_subscript0_share2_1 , x1x3x5x6_subscript0_share2_1 , x1x3x5x7_subscript0_share2_1 , x1x4x6x7_subscript0_share2_1 , x2x3x4x5_subscript0_share2_1 , x2x3x4x7_subscript0_share2_1 , x2x4x6x7_subscript0_share2_1 , x3x4x5x6_subscript0_share2_1 , x3x4x5x7_subscript0_share2_1 , x3x4x6x7_subscript0_share2_1 , x0x1x3x5_subscript0_share2_1 , x0x1x4x6_subscript0_share2_1 , x0x2x3x4_subscript0_share2_1 , x0x2x4x6_subscript0_share2_1 , x0x3x4x7_subscript0_share2_1 , x0x3x5x7_subscript0_share2_1 , x1x2x3x4_subscript0_share2_1 , x2x3x4x6_subscript0_share2_1 , x2x3x5x6_subscript0_share2_1 , x2x5x6x7_subscript0_share2_1 , x4x5x6x7_subscript0_share2_1 , x0x1x2x4_subscript0_share2_1 , x0x1x6x7_subscript0_share2_1 , x0x2x6x7_subscript0_share2_1 , x0x3x6x7_subscript0_share2_1 , x0x5x6x7_subscript0_share2_1 , x1x2x4x5_subscript0_share2_1 , x0x1x3x7_subscript0_share2_1 , x0x1x5x7_subscript0_share2_1 , x0x1x2x3x4_subscript0_share2_1 , x0x1x2x3x6_subscript0_share2_1 , x0x1x2x3x7_subscript0_share2_1 , x0x1x2x4x5_subscript0_share2_1 , x0x1x2x4x7_subscript0_share2_1 , x0x1x2x5x7_subscript0_share2_1 , x0x1x2x6x7_subscript0_share2_1 , x0x1x3x4x6_subscript0_share2_1 , x0x1x3x5x6_subscript0_share2_1 , x0x1x3x5x7_subscript0_share2_1 , x0x1x3x6x7_subscript0_share2_1 , x0x1x4x5x6_subscript0_share2_1 , x0x1x5x6x7_subscript0_share2_1 , x0x2x3x4x5_subscript0_share2_1 , x0x2x3x4x6_subscript0_share2_1 , x0x2x4x5x7_subscript0_share2_1 , x0x2x4x6x7_subscript0_share2_1 , x0x3x4x5x6_subscript0_share2_1 , x0x3x4x5x7_subscript0_share2_1 , x0x3x4x6x7_subscript0_share2_1 , x0x3x5x6x7_subscript0_share2_1 , x1x2x3x5x6_subscript0_share2_1 , x1x2x3x5x7_subscript0_share2_1 , x1x2x4x5x6_subscript0_share2_1 , x1x2x4x6x7_subscript0_share2_1 , x1x2x5x6x7_subscript0_share2_1 , x1x3x4x5x7_subscript0_share2_1 , x2x3x4x5x6_subscript0_share2_1 , x2x3x4x5x7_subscript0_share2_1 , x2x4x5x6x7_subscript0_share2_1 , x0x1x2x4x6_subscript0_share2_1 , x0x1x3x4x7_subscript0_share2_1 , x0x2x3x4x7_subscript0_share2_1 , x0x2x3x5x7_subscript0_share2_1 , x0x2x3x6x7_subscript0_share2_1 , x0x2x4x5x6_subscript0_share2_1 , x0x2x5x6x7_subscript0_share2_1 , x0x4x5x6x7_subscript0_share2_1 , x1x2x3x4x6_subscript0_share2_1 , x1x3x4x5x6_subscript0_share2_1 , x2x3x4x6x7_subscript0_share2_1 , x0x1x2x3x5_subscript0_share2_1 , x0x1x4x6x7_subscript0_share2_1 , x1x2x3x4x5_subscript0_share2_1 , x1x2x3x6x7_subscript0_share2_1 , x1x2x4x5x7_subscript0_share2_1 , x1x3x4x6x7_subscript0_share2_1 , x1x3x5x6x7_subscript0_share2_1 , x1x4x5x6x7_subscript0_share2_1 , x2x3x5x6x7_subscript0_share2_1 , x3x4x5x6x7_subscript0_share2_1 , x0x1x2x5x6_subscript0_share2_1 , x0x1x3x4x5_subscript0_share2_1 , x0x1x4x5x7_subscript0_share2_1 , x0x2x3x5x6_subscript0_share2_1 , x1x2x3x4x7_subscript0_share2_1 , x0x1x2x3x4x6_subscript0_share2_1 , x0x1x2x3x4x7_subscript0_share2_1 , x0x1x2x3x5x7_subscript0_share2_1 , x0x1x2x3x6x7_subscript0_share2_1 , x0x1x2x4x5x7_subscript0_share2_1 , x0x1x2x5x6x7_subscript0_share2_1 , x0x1x3x4x6x7_subscript0_share2_1 , x0x1x4x5x6x7_subscript0_share2_1 , x0x2x3x4x5x6_subscript0_share2_1 , x0x2x3x4x5x7_subscript0_share2_1 , x0x2x3x5x6x7_subscript0_share2_1 , x1x2x3x4x6x7_subscript0_share2_1 , x1x2x4x5x6x7_subscript0_share2_1 , x1x3x4x5x6x7_subscript0_share2_1 , x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x5x6_subscript0_share2_1 , x0x1x2x4x6x7_subscript0_share2_1 , x0x1x3x4x5x6_subscript0_share2_1 , x0x2x3x4x6x7_subscript0_share2_1 , x1x2x3x4x5x6_subscript0_share2_1 , x1x2x3x5x6x7_subscript0_share2_1 , x0x1x2x3x4x5_subscript0_share2_1 , x0x1x2x4x5x6_subscript0_share2_1 , x0x1x3x4x5x7_subscript0_share2_1 , x0x1x3x5x6x7_subscript0_share2_1 , x0x2x4x5x6x7_subscript0_share2_1 , x1x2x3x4x5x7_subscript0_share2_1 , x0x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x4x6x7_subscript0_share2_1 , x0x1x2x4x5x6x7_subscript0_share2_1 , x0x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x5x6x7_subscript0_share2_1 , x0x1x3x4x5x6x7_subscript0_share2_1 , x1x2x3x4x5x6x7_subscript0_share2_1 , x0x1x2x3x4x5x6_subscript0_share2_1 , x0x1x2x3x4x5x7_subscript0_share2_1 ;


wire  x0_share1 , x1_share1 , x2_share1 , x3_share1 , x4_share1 , x5_share1 , x6_share1 , x7_share1 ;

assign x0_share1 = input_share1[0] ^ rand_composable_bit[0] ;
assign x1_share1 = input_share1[1] ^ rand_composable_bit[1] ;
assign x2_share1 = input_share1[2] ^ rand_composable_bit[2] ;
assign x3_share1 = input_share1[3] ^ rand_composable_bit[3] ;
assign x4_share1 = input_share1[4] ^ rand_composable_bit[4] ;
assign x5_share1 = input_share1[5] ^ rand_composable_bit[5] ;
assign x6_share1 = input_share1[6] ^ rand_composable_bit[6] ;
assign x7_share1 = input_share1[7] ^ rand_composable_bit[7] ;




assign x0_subscript0_share1_1 = ( x0_share1 ) ^ rand_bit[1] ; 
assign x0_subscript0_share2_1 = rand_bit[1] ; 
assign x2_subscript0_share1_1 = ( x2_share1 ) ^ rand_bit[2] ; 
assign x2_subscript0_share2_1 = rand_bit[2] ; 
assign x3_subscript0_share1_1 = ( x3_share1 ) ^ rand_bit[3] ; 
assign x3_subscript0_share2_1 = rand_bit[3] ; 
assign x4_subscript0_share1_1 = ( x4_share1 ) ^ rand_bit[4] ; 
assign x4_subscript0_share2_1 = rand_bit[4] ; 
assign x6_subscript0_share1_1 = ( x6_share1 ) ^ rand_bit[5] ; 
assign x6_subscript0_share2_1 = rand_bit[5] ; 
assign x7_subscript0_share1_1 = ( x7_share1 ) ^ rand_bit[6] ; 
assign x7_subscript0_share2_1 = rand_bit[6] ; 
assign x1_subscript0_share1_1 = ( x1_share1 ) ^ rand_bit[7] ; 
assign x1_subscript0_share2_1 = rand_bit[7] ; 
assign x5_subscript0_share1_1 = ( x5_share1 ) ^ rand_bit[8] ; 
assign x5_subscript0_share2_1 = rand_bit[8] ; 
assign x0x1_subscript0_share1_1 = ( x0_share1 & x1_share1 ) ^ rand_bit[9] ; 
assign x0x1_subscript0_share2_1 = rand_bit[9] ; 
assign x0x4_subscript0_share1_1 = ( x0_share1 & x4_share1 ) ^ rand_bit[10] ; 
assign x0x4_subscript0_share2_1 = rand_bit[10] ; 
assign x0x5_subscript0_share1_1 = ( x0_share1 & x5_share1 ) ^ rand_bit[11] ; 
assign x0x5_subscript0_share2_1 = rand_bit[11] ; 
assign x0x6_subscript0_share1_1 = ( x0_share1 & x6_share1 ) ^ rand_bit[12] ; 
assign x0x6_subscript0_share2_1 = rand_bit[12] ; 
assign x1x2_subscript0_share1_1 = ( x1_share1 & x2_share1 ) ^ rand_bit[13] ; 
assign x1x2_subscript0_share2_1 = rand_bit[13] ; 
assign x1x3_subscript0_share1_1 = ( x1_share1 & x3_share1 ) ^ rand_bit[14] ; 
assign x1x3_subscript0_share2_1 = rand_bit[14] ; 
assign x1x4_subscript0_share1_1 = ( x1_share1 & x4_share1 ) ^ rand_bit[15] ; 
assign x1x4_subscript0_share2_1 = rand_bit[15] ; 
assign x1x6_subscript0_share1_1 = ( x1_share1 & x6_share1 ) ^ rand_bit[16] ; 
assign x1x6_subscript0_share2_1 = rand_bit[16] ; 
assign x2x3_subscript0_share1_1 = ( x2_share1 & x3_share1 ) ^ rand_bit[17] ; 
assign x2x3_subscript0_share2_1 = rand_bit[17] ; 
assign x2x4_subscript0_share1_1 = ( x2_share1 & x4_share1 ) ^ rand_bit[18] ; 
assign x2x4_subscript0_share2_1 = rand_bit[18] ; 
assign x2x6_subscript0_share1_1 = ( x2_share1 & x6_share1 ) ^ rand_bit[19] ; 
assign x2x6_subscript0_share2_1 = rand_bit[19] ; 
assign x2x7_subscript0_share1_1 = ( x2_share1 & x7_share1 ) ^ rand_bit[20] ; 
assign x2x7_subscript0_share2_1 = rand_bit[20] ; 
assign x4x6_subscript0_share1_1 = ( x4_share1 & x6_share1 ) ^ rand_bit[21] ; 
assign x4x6_subscript0_share2_1 = rand_bit[21] ; 
assign x5x6_subscript0_share1_1 = ( x5_share1 & x6_share1 ) ^ rand_bit[22] ; 
assign x5x6_subscript0_share2_1 = rand_bit[22] ; 
assign x5x7_subscript0_share1_1 = ( x5_share1 & x7_share1 ) ^ rand_bit[23] ; 
assign x5x7_subscript0_share2_1 = rand_bit[23] ; 
assign x6x7_subscript0_share1_1 = ( x6_share1 & x7_share1 ) ^ rand_bit[24] ; 
assign x6x7_subscript0_share2_1 = rand_bit[24] ; 
assign x0x2_subscript0_share1_1 = ( x0_share1 & x2_share1 ) ^ rand_bit[25] ; 
assign x0x2_subscript0_share2_1 = rand_bit[25] ; 
assign x0x3_subscript0_share1_1 = ( x0_share1 & x3_share1 ) ^ rand_bit[26] ; 
assign x0x3_subscript0_share2_1 = rand_bit[26] ; 
assign x0x7_subscript0_share1_1 = ( x0_share1 & x7_share1 ) ^ rand_bit[27] ; 
assign x0x7_subscript0_share2_1 = rand_bit[27] ; 
assign x1x7_subscript0_share1_1 = ( x1_share1 & x7_share1 ) ^ rand_bit[28] ; 
assign x1x7_subscript0_share2_1 = rand_bit[28] ; 
assign x3x7_subscript0_share1_1 = ( x3_share1 & x7_share1 ) ^ rand_bit[29] ; 
assign x3x7_subscript0_share2_1 = rand_bit[29] ; 
assign x4x5_subscript0_share1_1 = ( x4_share1 & x5_share1 ) ^ rand_bit[30] ; 
assign x4x5_subscript0_share2_1 = rand_bit[30] ; 
assign x3x4_subscript0_share1_1 = ( x3_share1 & x4_share1 ) ^ rand_bit[31] ; 
assign x3x4_subscript0_share2_1 = rand_bit[31] ; 
assign x4x7_subscript0_share1_1 = ( x4_share1 & x7_share1 ) ^ rand_bit[32] ; 
assign x4x7_subscript0_share2_1 = rand_bit[32] ; 
assign x3x6_subscript0_share1_1 = ( x3_share1 & x6_share1 ) ^ rand_bit[33] ; 
assign x3x6_subscript0_share2_1 = rand_bit[33] ; 
assign x1x5_subscript0_share1_1 = ( x1_share1 & x5_share1 ) ^ rand_bit[34] ; 
assign x1x5_subscript0_share2_1 = rand_bit[34] ; 
assign x2x5_subscript0_share1_1 = ( x2_share1 & x5_share1 ) ^ rand_bit[35] ; 
assign x2x5_subscript0_share2_1 = rand_bit[35] ; 
assign x3x5_subscript0_share1_1 = ( x3_share1 & x5_share1 ) ^ rand_bit[36] ; 
assign x3x5_subscript0_share2_1 = rand_bit[36] ; 
assign x0x1x4_subscript0_share1_1 = ( x0_share1 & x1_share1 & x4_share1 ) ^ rand_bit[37] ; 
assign x0x1x4_subscript0_share2_1 = rand_bit[37] ; 
assign x0x1x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x6_share1 ) ^ rand_bit[38] ; 
assign x0x1x6_subscript0_share2_1 = rand_bit[38] ; 
assign x0x1x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x7_share1 ) ^ rand_bit[39] ; 
assign x0x1x7_subscript0_share2_1 = rand_bit[39] ; 
assign x0x2x4_subscript0_share1_1 = ( x0_share1 & x2_share1 & x4_share1 ) ^ rand_bit[40] ; 
assign x0x2x4_subscript0_share2_1 = rand_bit[40] ; 
assign x0x2x5_subscript0_share1_1 = ( x0_share1 & x2_share1 & x5_share1 ) ^ rand_bit[41] ; 
assign x0x2x5_subscript0_share2_1 = rand_bit[41] ; 
assign x0x2x6_subscript0_share1_1 = ( x0_share1 & x2_share1 & x6_share1 ) ^ rand_bit[42] ; 
assign x0x2x6_subscript0_share2_1 = rand_bit[42] ; 
assign x0x2x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x7_share1 ) ^ rand_bit[43] ; 
assign x0x2x7_subscript0_share2_1 = rand_bit[43] ; 
assign x0x3x4_subscript0_share1_1 = ( x0_share1 & x3_share1 & x4_share1 ) ^ rand_bit[44] ; 
assign x0x3x4_subscript0_share2_1 = rand_bit[44] ; 
assign x0x3x5_subscript0_share1_1 = ( x0_share1 & x3_share1 & x5_share1 ) ^ rand_bit[45] ; 
assign x0x3x5_subscript0_share2_1 = rand_bit[45] ; 
assign x0x3x6_subscript0_share1_1 = ( x0_share1 & x3_share1 & x6_share1 ) ^ rand_bit[46] ; 
assign x0x3x6_subscript0_share2_1 = rand_bit[46] ; 
assign x0x4x6_subscript0_share1_1 = ( x0_share1 & x4_share1 & x6_share1 ) ^ rand_bit[47] ; 
assign x0x4x6_subscript0_share2_1 = rand_bit[47] ; 
assign x0x4x7_subscript0_share1_1 = ( x0_share1 & x4_share1 & x7_share1 ) ^ rand_bit[48] ; 
assign x0x4x7_subscript0_share2_1 = rand_bit[48] ; 
assign x1x2x3_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 ) ^ rand_bit[49] ; 
assign x1x2x3_subscript0_share2_1 = rand_bit[49] ; 
assign x1x2x4_subscript0_share1_1 = ( x1_share1 & x2_share1 & x4_share1 ) ^ rand_bit[50] ; 
assign x1x2x4_subscript0_share2_1 = rand_bit[50] ; 
assign x1x2x6_subscript0_share1_1 = ( x1_share1 & x2_share1 & x6_share1 ) ^ rand_bit[51] ; 
assign x1x2x6_subscript0_share2_1 = rand_bit[51] ; 
assign x1x3x4_subscript0_share1_1 = ( x1_share1 & x3_share1 & x4_share1 ) ^ rand_bit[52] ; 
assign x1x3x4_subscript0_share2_1 = rand_bit[52] ; 
assign x1x3x7_subscript0_share1_1 = ( x1_share1 & x3_share1 & x7_share1 ) ^ rand_bit[53] ; 
assign x1x3x7_subscript0_share2_1 = rand_bit[53] ; 
assign x1x4x6_subscript0_share1_1 = ( x1_share1 & x4_share1 & x6_share1 ) ^ rand_bit[54] ; 
assign x1x4x6_subscript0_share2_1 = rand_bit[54] ; 
assign x1x5x6_subscript0_share1_1 = ( x1_share1 & x5_share1 & x6_share1 ) ^ rand_bit[55] ; 
assign x1x5x6_subscript0_share2_1 = rand_bit[55] ; 
assign x2x3x5_subscript0_share1_1 = ( x2_share1 & x3_share1 & x5_share1 ) ^ rand_bit[56] ; 
assign x2x3x5_subscript0_share2_1 = rand_bit[56] ; 
assign x2x3x7_subscript0_share1_1 = ( x2_share1 & x3_share1 & x7_share1 ) ^ rand_bit[57] ; 
assign x2x3x7_subscript0_share2_1 = rand_bit[57] ; 
assign x2x4x7_subscript0_share1_1 = ( x2_share1 & x4_share1 & x7_share1 ) ^ rand_bit[58] ; 
assign x2x4x7_subscript0_share2_1 = rand_bit[58] ; 
assign x2x5x6_subscript0_share1_1 = ( x2_share1 & x5_share1 & x6_share1 ) ^ rand_bit[59] ; 
assign x2x5x6_subscript0_share2_1 = rand_bit[59] ; 
assign x2x5x7_subscript0_share1_1 = ( x2_share1 & x5_share1 & x7_share1 ) ^ rand_bit[60] ; 
assign x2x5x7_subscript0_share2_1 = rand_bit[60] ; 
assign x2x6x7_subscript0_share1_1 = ( x2_share1 & x6_share1 & x7_share1 ) ^ rand_bit[61] ; 
assign x2x6x7_subscript0_share2_1 = rand_bit[61] ; 
assign x3x4x7_subscript0_share1_1 = ( x3_share1 & x4_share1 & x7_share1 ) ^ rand_bit[62] ; 
assign x3x4x7_subscript0_share2_1 = rand_bit[62] ; 
assign x3x5x7_subscript0_share1_1 = ( x3_share1 & x5_share1 & x7_share1 ) ^ rand_bit[63] ; 
assign x3x5x7_subscript0_share2_1 = rand_bit[63] ; 
assign x3x6x7_subscript0_share1_1 = ( x3_share1 & x6_share1 & x7_share1 ) ^ rand_bit[64] ; 
assign x3x6x7_subscript0_share2_1 = rand_bit[64] ; 
assign x4x5x6_subscript0_share1_1 = ( x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[65] ; 
assign x4x5x6_subscript0_share2_1 = rand_bit[65] ; 
assign x5x6x7_subscript0_share1_1 = ( x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[66] ; 
assign x5x6x7_subscript0_share2_1 = rand_bit[66] ; 
assign x0x1x3_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 ) ^ rand_bit[67] ; 
assign x0x1x3_subscript0_share2_1 = rand_bit[67] ; 
assign x0x2x3_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 ) ^ rand_bit[68] ; 
assign x0x2x3_subscript0_share2_1 = rand_bit[68] ; 
assign x0x4x5_subscript0_share1_1 = ( x0_share1 & x4_share1 & x5_share1 ) ^ rand_bit[69] ; 
assign x0x4x5_subscript0_share2_1 = rand_bit[69] ; 
assign x0x5x7_subscript0_share1_1 = ( x0_share1 & x5_share1 & x7_share1 ) ^ rand_bit[70] ; 
assign x0x5x7_subscript0_share2_1 = rand_bit[70] ; 
assign x0x6x7_subscript0_share1_1 = ( x0_share1 & x6_share1 & x7_share1 ) ^ rand_bit[71] ; 
assign x0x6x7_subscript0_share2_1 = rand_bit[71] ; 
assign x1x3x5_subscript0_share1_1 = ( x1_share1 & x3_share1 & x5_share1 ) ^ rand_bit[72] ; 
assign x1x3x5_subscript0_share2_1 = rand_bit[72] ; 
assign x1x3x6_subscript0_share1_1 = ( x1_share1 & x3_share1 & x6_share1 ) ^ rand_bit[73] ; 
assign x1x3x6_subscript0_share2_1 = rand_bit[73] ; 
assign x1x4x7_subscript0_share1_1 = ( x1_share1 & x4_share1 & x7_share1 ) ^ rand_bit[74] ; 
assign x1x4x7_subscript0_share2_1 = rand_bit[74] ; 
assign x2x3x4_subscript0_share1_1 = ( x2_share1 & x3_share1 & x4_share1 ) ^ rand_bit[75] ; 
assign x2x3x4_subscript0_share2_1 = rand_bit[75] ; 
assign x2x3x6_subscript0_share1_1 = ( x2_share1 & x3_share1 & x6_share1 ) ^ rand_bit[76] ; 
assign x2x3x6_subscript0_share2_1 = rand_bit[76] ; 
assign x3x4x6_subscript0_share1_1 = ( x3_share1 & x4_share1 & x6_share1 ) ^ rand_bit[77] ; 
assign x3x4x6_subscript0_share2_1 = rand_bit[77] ; 
assign x3x5x6_subscript0_share1_1 = ( x3_share1 & x5_share1 & x6_share1 ) ^ rand_bit[78] ; 
assign x3x5x6_subscript0_share2_1 = rand_bit[78] ; 
assign x0x1x5_subscript0_share1_1 = ( x0_share1 & x1_share1 & x5_share1 ) ^ rand_bit[79] ; 
assign x0x1x5_subscript0_share2_1 = rand_bit[79] ; 
assign x0x3x7_subscript0_share1_1 = ( x0_share1 & x3_share1 & x7_share1 ) ^ rand_bit[80] ; 
assign x0x3x7_subscript0_share2_1 = rand_bit[80] ; 
assign x1x2x5_subscript0_share1_1 = ( x1_share1 & x2_share1 & x5_share1 ) ^ rand_bit[81] ; 
assign x1x2x5_subscript0_share2_1 = rand_bit[81] ; 
assign x1x2x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x7_share1 ) ^ rand_bit[82] ; 
assign x1x2x7_subscript0_share2_1 = rand_bit[82] ; 
assign x1x4x5_subscript0_share1_1 = ( x1_share1 & x4_share1 & x5_share1 ) ^ rand_bit[83] ; 
assign x1x4x5_subscript0_share2_1 = rand_bit[83] ; 
assign x1x5x7_subscript0_share1_1 = ( x1_share1 & x5_share1 & x7_share1 ) ^ rand_bit[84] ; 
assign x1x5x7_subscript0_share2_1 = rand_bit[84] ; 
assign x2x4x5_subscript0_share1_1 = ( x2_share1 & x4_share1 & x5_share1 ) ^ rand_bit[85] ; 
assign x2x4x5_subscript0_share2_1 = rand_bit[85] ; 
assign x3x4x5_subscript0_share1_1 = ( x3_share1 & x4_share1 & x5_share1 ) ^ rand_bit[86] ; 
assign x3x4x5_subscript0_share2_1 = rand_bit[86] ; 
assign x4x6x7_subscript0_share1_1 = ( x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[87] ; 
assign x4x6x7_subscript0_share2_1 = rand_bit[87] ; 
assign x1x6x7_subscript0_share1_1 = ( x1_share1 & x6_share1 & x7_share1 ) ^ rand_bit[88] ; 
assign x1x6x7_subscript0_share2_1 = rand_bit[88] ; 
assign x4x5x7_subscript0_share1_1 = ( x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[89] ; 
assign x4x5x7_subscript0_share2_1 = rand_bit[89] ; 
assign x0x1x2_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 ) ^ rand_bit[90] ; 
assign x0x1x2_subscript0_share2_1 = rand_bit[90] ; 
assign x0x5x6_subscript0_share1_1 = ( x0_share1 & x5_share1 & x6_share1 ) ^ rand_bit[91] ; 
assign x0x5x6_subscript0_share2_1 = rand_bit[91] ; 
assign x2x4x6_subscript0_share1_1 = ( x2_share1 & x4_share1 & x6_share1 ) ^ rand_bit[92] ; 
assign x2x4x6_subscript0_share2_1 = rand_bit[92] ; 
assign x0x1x2x3_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 ) ^ rand_bit[93] ; 
assign x0x1x2x3_subscript0_share2_1 = rand_bit[93] ; 
assign x0x1x2x5_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x5_share1 ) ^ rand_bit[94] ; 
assign x0x1x2x5_subscript0_share2_1 = rand_bit[94] ; 
assign x0x1x2x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x6_share1 ) ^ rand_bit[95] ; 
assign x0x1x2x6_subscript0_share2_1 = rand_bit[95] ; 
assign x0x1x2x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x7_share1 ) ^ rand_bit[96] ; 
assign x0x1x2x7_subscript0_share2_1 = rand_bit[96] ; 
assign x0x1x4x5_subscript0_share1_1 = ( x0_share1 & x1_share1 & x4_share1 & x5_share1 ) ^ rand_bit[97] ; 
assign x0x1x4x5_subscript0_share2_1 = rand_bit[97] ; 
assign x0x1x4x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x4_share1 & x7_share1 ) ^ rand_bit[98] ; 
assign x0x1x4x7_subscript0_share2_1 = rand_bit[98] ; 
assign x0x2x3x5_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x5_share1 ) ^ rand_bit[99] ; 
assign x0x2x3x5_subscript0_share2_1 = rand_bit[99] ; 
assign x0x2x3x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x7_share1 ) ^ rand_bit[100] ; 
assign x0x2x3x7_subscript0_share2_1 = rand_bit[100] ; 
assign x0x2x4x5_subscript0_share1_1 = ( x0_share1 & x2_share1 & x4_share1 & x5_share1 ) ^ rand_bit[101] ; 
assign x0x2x4x5_subscript0_share2_1 = rand_bit[101] ; 
assign x0x2x4x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x4_share1 & x7_share1 ) ^ rand_bit[102] ; 
assign x0x2x4x7_subscript0_share2_1 = rand_bit[102] ; 
assign x0x2x5x6_subscript0_share1_1 = ( x0_share1 & x2_share1 & x5_share1 & x6_share1 ) ^ rand_bit[103] ; 
assign x0x2x5x6_subscript0_share2_1 = rand_bit[103] ; 
assign x0x2x5x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x5_share1 & x7_share1 ) ^ rand_bit[104] ; 
assign x0x2x5x7_subscript0_share2_1 = rand_bit[104] ; 
assign x0x3x4x6_subscript0_share1_1 = ( x0_share1 & x3_share1 & x4_share1 & x6_share1 ) ^ rand_bit[105] ; 
assign x0x3x4x6_subscript0_share2_1 = rand_bit[105] ; 
assign x0x3x5x6_subscript0_share1_1 = ( x0_share1 & x3_share1 & x5_share1 & x6_share1 ) ^ rand_bit[106] ; 
assign x0x3x5x6_subscript0_share2_1 = rand_bit[106] ; 
assign x0x4x5x6_subscript0_share1_1 = ( x0_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[107] ; 
assign x0x4x5x6_subscript0_share2_1 = rand_bit[107] ; 
assign x0x4x5x7_subscript0_share1_1 = ( x0_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[108] ; 
assign x0x4x5x7_subscript0_share2_1 = rand_bit[108] ; 
assign x0x4x6x7_subscript0_share1_1 = ( x0_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[109] ; 
assign x0x4x6x7_subscript0_share2_1 = rand_bit[109] ; 
assign x1x2x3x5_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x5_share1 ) ^ rand_bit[110] ; 
assign x1x2x3x5_subscript0_share2_1 = rand_bit[110] ; 
assign x1x2x3x6_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x6_share1 ) ^ rand_bit[111] ; 
assign x1x2x3x6_subscript0_share2_1 = rand_bit[111] ; 
assign x1x2x3x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x7_share1 ) ^ rand_bit[112] ; 
assign x1x2x3x7_subscript0_share2_1 = rand_bit[112] ; 
assign x1x2x4x6_subscript0_share1_1 = ( x1_share1 & x2_share1 & x4_share1 & x6_share1 ) ^ rand_bit[113] ; 
assign x1x2x4x6_subscript0_share2_1 = rand_bit[113] ; 
assign x1x2x4x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x4_share1 & x7_share1 ) ^ rand_bit[114] ; 
assign x1x2x4x7_subscript0_share2_1 = rand_bit[114] ; 
assign x1x2x6x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x6_share1 & x7_share1 ) ^ rand_bit[115] ; 
assign x1x2x6x7_subscript0_share2_1 = rand_bit[115] ; 
assign x1x3x4x6_subscript0_share1_1 = ( x1_share1 & x3_share1 & x4_share1 & x6_share1 ) ^ rand_bit[116] ; 
assign x1x3x4x6_subscript0_share2_1 = rand_bit[116] ; 
assign x1x3x6x7_subscript0_share1_1 = ( x1_share1 & x3_share1 & x6_share1 & x7_share1 ) ^ rand_bit[117] ; 
assign x1x3x6x7_subscript0_share2_1 = rand_bit[117] ; 
assign x1x4x5x6_subscript0_share1_1 = ( x1_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[118] ; 
assign x1x4x5x6_subscript0_share2_1 = rand_bit[118] ; 
assign x1x4x5x7_subscript0_share1_1 = ( x1_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[119] ; 
assign x1x4x5x7_subscript0_share2_1 = rand_bit[119] ; 
assign x1x5x6x7_subscript0_share1_1 = ( x1_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[120] ; 
assign x1x5x6x7_subscript0_share2_1 = rand_bit[120] ; 
assign x2x3x5x7_subscript0_share1_1 = ( x2_share1 & x3_share1 & x5_share1 & x7_share1 ) ^ rand_bit[121] ; 
assign x2x3x5x7_subscript0_share2_1 = rand_bit[121] ; 
assign x2x3x6x7_subscript0_share1_1 = ( x2_share1 & x3_share1 & x6_share1 & x7_share1 ) ^ rand_bit[122] ; 
assign x2x3x6x7_subscript0_share2_1 = rand_bit[122] ; 
assign x2x4x5x6_subscript0_share1_1 = ( x2_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[123] ; 
assign x2x4x5x6_subscript0_share2_1 = rand_bit[123] ; 
assign x2x4x5x7_subscript0_share1_1 = ( x2_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[124] ; 
assign x2x4x5x7_subscript0_share2_1 = rand_bit[124] ; 
assign x3x5x6x7_subscript0_share1_1 = ( x3_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[125] ; 
assign x3x5x6x7_subscript0_share2_1 = rand_bit[125] ; 
assign x0x1x3x4_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x4_share1 ) ^ rand_bit[126] ; 
assign x0x1x3x4_subscript0_share2_1 = rand_bit[126] ; 
assign x0x1x3x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x6_share1 ) ^ rand_bit[127] ; 
assign x0x1x3x6_subscript0_share2_1 = rand_bit[127] ; 
assign x0x1x5x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x5_share1 & x6_share1 ) ^ rand_bit[128] ; 
assign x0x1x5x6_subscript0_share2_1 = rand_bit[128] ; 
assign x0x2x3x6_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x6_share1 ) ^ rand_bit[129] ; 
assign x0x2x3x6_subscript0_share2_1 = rand_bit[129] ; 
assign x0x3x4x5_subscript0_share1_1 = ( x0_share1 & x3_share1 & x4_share1 & x5_share1 ) ^ rand_bit[130] ; 
assign x0x3x4x5_subscript0_share2_1 = rand_bit[130] ; 
assign x1x2x5x6_subscript0_share1_1 = ( x1_share1 & x2_share1 & x5_share1 & x6_share1 ) ^ rand_bit[131] ; 
assign x1x2x5x6_subscript0_share2_1 = rand_bit[131] ; 
assign x1x2x5x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x5_share1 & x7_share1 ) ^ rand_bit[132] ; 
assign x1x2x5x7_subscript0_share2_1 = rand_bit[132] ; 
assign x1x3x4x5_subscript0_share1_1 = ( x1_share1 & x3_share1 & x4_share1 & x5_share1 ) ^ rand_bit[133] ; 
assign x1x3x4x5_subscript0_share2_1 = rand_bit[133] ; 
assign x1x3x4x7_subscript0_share1_1 = ( x1_share1 & x3_share1 & x4_share1 & x7_share1 ) ^ rand_bit[134] ; 
assign x1x3x4x7_subscript0_share2_1 = rand_bit[134] ; 
assign x1x3x5x6_subscript0_share1_1 = ( x1_share1 & x3_share1 & x5_share1 & x6_share1 ) ^ rand_bit[135] ; 
assign x1x3x5x6_subscript0_share2_1 = rand_bit[135] ; 
assign x1x3x5x7_subscript0_share1_1 = ( x1_share1 & x3_share1 & x5_share1 & x7_share1 ) ^ rand_bit[136] ; 
assign x1x3x5x7_subscript0_share2_1 = rand_bit[136] ; 
assign x1x4x6x7_subscript0_share1_1 = ( x1_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[137] ; 
assign x1x4x6x7_subscript0_share2_1 = rand_bit[137] ; 
assign x2x3x4x5_subscript0_share1_1 = ( x2_share1 & x3_share1 & x4_share1 & x5_share1 ) ^ rand_bit[138] ; 
assign x2x3x4x5_subscript0_share2_1 = rand_bit[138] ; 
assign x2x3x4x7_subscript0_share1_1 = ( x2_share1 & x3_share1 & x4_share1 & x7_share1 ) ^ rand_bit[139] ; 
assign x2x3x4x7_subscript0_share2_1 = rand_bit[139] ; 
assign x2x4x6x7_subscript0_share1_1 = ( x2_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[140] ; 
assign x2x4x6x7_subscript0_share2_1 = rand_bit[140] ; 
assign x3x4x5x6_subscript0_share1_1 = ( x3_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[141] ; 
assign x3x4x5x6_subscript0_share2_1 = rand_bit[141] ; 
assign x3x4x5x7_subscript0_share1_1 = ( x3_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[142] ; 
assign x3x4x5x7_subscript0_share2_1 = rand_bit[142] ; 
assign x3x4x6x7_subscript0_share1_1 = ( x3_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[143] ; 
assign x3x4x6x7_subscript0_share2_1 = rand_bit[143] ; 
assign x0x1x3x5_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x5_share1 ) ^ rand_bit[144] ; 
assign x0x1x3x5_subscript0_share2_1 = rand_bit[144] ; 
assign x0x1x4x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x4_share1 & x6_share1 ) ^ rand_bit[145] ; 
assign x0x1x4x6_subscript0_share2_1 = rand_bit[145] ; 
assign x0x2x3x4_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x4_share1 ) ^ rand_bit[146] ; 
assign x0x2x3x4_subscript0_share2_1 = rand_bit[146] ; 
assign x0x2x4x6_subscript0_share1_1 = ( x0_share1 & x2_share1 & x4_share1 & x6_share1 ) ^ rand_bit[147] ; 
assign x0x2x4x6_subscript0_share2_1 = rand_bit[147] ; 
assign x0x3x4x7_subscript0_share1_1 = ( x0_share1 & x3_share1 & x4_share1 & x7_share1 ) ^ rand_bit[148] ; 
assign x0x3x4x7_subscript0_share2_1 = rand_bit[148] ; 
assign x0x3x5x7_subscript0_share1_1 = ( x0_share1 & x3_share1 & x5_share1 & x7_share1 ) ^ rand_bit[149] ; 
assign x0x3x5x7_subscript0_share2_1 = rand_bit[149] ; 
assign x1x2x3x4_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x4_share1 ) ^ rand_bit[150] ; 
assign x1x2x3x4_subscript0_share2_1 = rand_bit[150] ; 
assign x2x3x4x6_subscript0_share1_1 = ( x2_share1 & x3_share1 & x4_share1 & x6_share1 ) ^ rand_bit[151] ; 
assign x2x3x4x6_subscript0_share2_1 = rand_bit[151] ; 
assign x2x3x5x6_subscript0_share1_1 = ( x2_share1 & x3_share1 & x5_share1 & x6_share1 ) ^ rand_bit[152] ; 
assign x2x3x5x6_subscript0_share2_1 = rand_bit[152] ; 
assign x2x5x6x7_subscript0_share1_1 = ( x2_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[153] ; 
assign x2x5x6x7_subscript0_share2_1 = rand_bit[153] ; 
assign x4x5x6x7_subscript0_share1_1 = ( x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[154] ; 
assign x4x5x6x7_subscript0_share2_1 = rand_bit[154] ; 
assign x0x1x2x4_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x4_share1 ) ^ rand_bit[155] ; 
assign x0x1x2x4_subscript0_share2_1 = rand_bit[155] ; 
assign x0x1x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x6_share1 & x7_share1 ) ^ rand_bit[156] ; 
assign x0x1x6x7_subscript0_share2_1 = rand_bit[156] ; 
assign x0x2x6x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x6_share1 & x7_share1 ) ^ rand_bit[157] ; 
assign x0x2x6x7_subscript0_share2_1 = rand_bit[157] ; 
assign x0x3x6x7_subscript0_share1_1 = ( x0_share1 & x3_share1 & x6_share1 & x7_share1 ) ^ rand_bit[158] ; 
assign x0x3x6x7_subscript0_share2_1 = rand_bit[158] ; 
assign x0x5x6x7_subscript0_share1_1 = ( x0_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[159] ; 
assign x0x5x6x7_subscript0_share2_1 = rand_bit[159] ; 
assign x1x2x4x5_subscript0_share1_1 = ( x1_share1 & x2_share1 & x4_share1 & x5_share1 ) ^ rand_bit[160] ; 
assign x1x2x4x5_subscript0_share2_1 = rand_bit[160] ; 
assign x0x1x3x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x7_share1 ) ^ rand_bit[161] ; 
assign x0x1x3x7_subscript0_share2_1 = rand_bit[161] ; 
assign x0x1x5x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x5_share1 & x7_share1 ) ^ rand_bit[162] ; 
assign x0x1x5x7_subscript0_share2_1 = rand_bit[162] ; 
assign x0x1x2x3x4_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x4_share1 ) ^ rand_bit[163] ; 
assign x0x1x2x3x4_subscript0_share2_1 = rand_bit[163] ; 
assign x0x1x2x3x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x6_share1 ) ^ rand_bit[164] ; 
assign x0x1x2x3x6_subscript0_share2_1 = rand_bit[164] ; 
assign x0x1x2x3x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x7_share1 ) ^ rand_bit[165] ; 
assign x0x1x2x3x7_subscript0_share2_1 = rand_bit[165] ; 
assign x0x1x2x4x5_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x4_share1 & x5_share1 ) ^ rand_bit[166] ; 
assign x0x1x2x4x5_subscript0_share2_1 = rand_bit[166] ; 
assign x0x1x2x4x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x4_share1 & x7_share1 ) ^ rand_bit[167] ; 
assign x0x1x2x4x7_subscript0_share2_1 = rand_bit[167] ; 
assign x0x1x2x5x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x5_share1 & x7_share1 ) ^ rand_bit[168] ; 
assign x0x1x2x5x7_subscript0_share2_1 = rand_bit[168] ; 
assign x0x1x2x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x6_share1 & x7_share1 ) ^ rand_bit[169] ; 
assign x0x1x2x6x7_subscript0_share2_1 = rand_bit[169] ; 
assign x0x1x3x4x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x4_share1 & x6_share1 ) ^ rand_bit[170] ; 
assign x0x1x3x4x6_subscript0_share2_1 = rand_bit[170] ; 
assign x0x1x3x5x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x5_share1 & x6_share1 ) ^ rand_bit[171] ; 
assign x0x1x3x5x6_subscript0_share2_1 = rand_bit[171] ; 
assign x0x1x3x5x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x5_share1 & x7_share1 ) ^ rand_bit[172] ; 
assign x0x1x3x5x7_subscript0_share2_1 = rand_bit[172] ; 
assign x0x1x3x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x6_share1 & x7_share1 ) ^ rand_bit[173] ; 
assign x0x1x3x6x7_subscript0_share2_1 = rand_bit[173] ; 
assign x0x1x4x5x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[174] ; 
assign x0x1x4x5x6_subscript0_share2_1 = rand_bit[174] ; 
assign x0x1x5x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[175] ; 
assign x0x1x5x6x7_subscript0_share2_1 = rand_bit[175] ; 
assign x0x2x3x4x5_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 ) ^ rand_bit[176] ; 
assign x0x2x3x4x5_subscript0_share2_1 = rand_bit[176] ; 
assign x0x2x3x4x6_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x4_share1 & x6_share1 ) ^ rand_bit[177] ; 
assign x0x2x3x4x6_subscript0_share2_1 = rand_bit[177] ; 
assign x0x2x4x5x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[178] ; 
assign x0x2x4x5x7_subscript0_share2_1 = rand_bit[178] ; 
assign x0x2x4x6x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[179] ; 
assign x0x2x4x6x7_subscript0_share2_1 = rand_bit[179] ; 
assign x0x3x4x5x6_subscript0_share1_1 = ( x0_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[180] ; 
assign x0x3x4x5x6_subscript0_share2_1 = rand_bit[180] ; 
assign x0x3x4x5x7_subscript0_share1_1 = ( x0_share1 & x3_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[181] ; 
assign x0x3x4x5x7_subscript0_share2_1 = rand_bit[181] ; 
assign x0x3x4x6x7_subscript0_share1_1 = ( x0_share1 & x3_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[182] ; 
assign x0x3x4x6x7_subscript0_share2_1 = rand_bit[182] ; 
assign x0x3x5x6x7_subscript0_share1_1 = ( x0_share1 & x3_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[183] ; 
assign x0x3x5x6x7_subscript0_share2_1 = rand_bit[183] ; 
assign x1x2x3x5x6_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x5_share1 & x6_share1 ) ^ rand_bit[184] ; 
assign x1x2x3x5x6_subscript0_share2_1 = rand_bit[184] ; 
assign x1x2x3x5x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x5_share1 & x7_share1 ) ^ rand_bit[185] ; 
assign x1x2x3x5x7_subscript0_share2_1 = rand_bit[185] ; 
assign x1x2x4x5x6_subscript0_share1_1 = ( x1_share1 & x2_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[186] ; 
assign x1x2x4x5x6_subscript0_share2_1 = rand_bit[186] ; 
assign x1x2x4x6x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[187] ; 
assign x1x2x4x6x7_subscript0_share2_1 = rand_bit[187] ; 
assign x1x2x5x6x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[188] ; 
assign x1x2x5x6x7_subscript0_share2_1 = rand_bit[188] ; 
assign x1x3x4x5x7_subscript0_share1_1 = ( x1_share1 & x3_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[189] ; 
assign x1x3x4x5x7_subscript0_share2_1 = rand_bit[189] ; 
assign x2x3x4x5x6_subscript0_share1_1 = ( x2_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[190] ; 
assign x2x3x4x5x6_subscript0_share2_1 = rand_bit[190] ; 
assign x2x3x4x5x7_subscript0_share1_1 = ( x2_share1 & x3_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[191] ; 
assign x2x3x4x5x7_subscript0_share2_1 = rand_bit[191] ; 
assign x2x4x5x6x7_subscript0_share1_1 = ( x2_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[192] ; 
assign x2x4x5x6x7_subscript0_share2_1 = rand_bit[192] ; 
assign x0x1x2x4x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x4_share1 & x6_share1 ) ^ rand_bit[193] ; 
assign x0x1x2x4x6_subscript0_share2_1 = rand_bit[193] ; 
assign x0x1x3x4x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x4_share1 & x7_share1 ) ^ rand_bit[194] ; 
assign x0x1x3x4x7_subscript0_share2_1 = rand_bit[194] ; 
assign x0x2x3x4x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x4_share1 & x7_share1 ) ^ rand_bit[195] ; 
assign x0x2x3x4x7_subscript0_share2_1 = rand_bit[195] ; 
assign x0x2x3x5x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x5_share1 & x7_share1 ) ^ rand_bit[196] ; 
assign x0x2x3x5x7_subscript0_share2_1 = rand_bit[196] ; 
assign x0x2x3x6x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x6_share1 & x7_share1 ) ^ rand_bit[197] ; 
assign x0x2x3x6x7_subscript0_share2_1 = rand_bit[197] ; 
assign x0x2x4x5x6_subscript0_share1_1 = ( x0_share1 & x2_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[198] ; 
assign x0x2x4x5x6_subscript0_share2_1 = rand_bit[198] ; 
assign x0x2x5x6x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[199] ; 
assign x0x2x5x6x7_subscript0_share2_1 = rand_bit[199] ; 
assign x0x4x5x6x7_subscript0_share1_1 = ( x0_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[200] ; 
assign x0x4x5x6x7_subscript0_share2_1 = rand_bit[200] ; 
assign x1x2x3x4x6_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x4_share1 & x6_share1 ) ^ rand_bit[201] ; 
assign x1x2x3x4x6_subscript0_share2_1 = rand_bit[201] ; 
assign x1x3x4x5x6_subscript0_share1_1 = ( x1_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[202] ; 
assign x1x3x4x5x6_subscript0_share2_1 = rand_bit[202] ; 
assign x2x3x4x6x7_subscript0_share1_1 = ( x2_share1 & x3_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[203] ; 
assign x2x3x4x6x7_subscript0_share2_1 = rand_bit[203] ; 
assign x0x1x2x3x5_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x5_share1 ) ^ rand_bit[204] ; 
assign x0x1x2x3x5_subscript0_share2_1 = rand_bit[204] ; 
assign x0x1x4x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[205] ; 
assign x0x1x4x6x7_subscript0_share2_1 = rand_bit[205] ; 
assign x1x2x3x4x5_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 ) ^ rand_bit[206] ; 
assign x1x2x3x4x5_subscript0_share2_1 = rand_bit[206] ; 
assign x1x2x3x6x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x6_share1 & x7_share1 ) ^ rand_bit[207] ; 
assign x1x2x3x6x7_subscript0_share2_1 = rand_bit[207] ; 
assign x1x2x4x5x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[208] ; 
assign x1x2x4x5x7_subscript0_share2_1 = rand_bit[208] ; 
assign x1x3x4x6x7_subscript0_share1_1 = ( x1_share1 & x3_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[209] ; 
assign x1x3x4x6x7_subscript0_share2_1 = rand_bit[209] ; 
assign x1x3x5x6x7_subscript0_share1_1 = ( x1_share1 & x3_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[210] ; 
assign x1x3x5x6x7_subscript0_share2_1 = rand_bit[210] ; 
assign x1x4x5x6x7_subscript0_share1_1 = ( x1_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[211] ; 
assign x1x4x5x6x7_subscript0_share2_1 = rand_bit[211] ; 
assign x2x3x5x6x7_subscript0_share1_1 = ( x2_share1 & x3_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[212] ; 
assign x2x3x5x6x7_subscript0_share2_1 = rand_bit[212] ; 
assign x3x4x5x6x7_subscript0_share1_1 = ( x3_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[213] ; 
assign x3x4x5x6x7_subscript0_share2_1 = rand_bit[213] ; 
assign x0x1x2x5x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x5_share1 & x6_share1 ) ^ rand_bit[214] ; 
assign x0x1x2x5x6_subscript0_share2_1 = rand_bit[214] ; 
assign x0x1x3x4x5_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x4_share1 & x5_share1 ) ^ rand_bit[215] ; 
assign x0x1x3x4x5_subscript0_share2_1 = rand_bit[215] ; 
assign x0x1x4x5x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[216] ; 
assign x0x1x4x5x7_subscript0_share2_1 = rand_bit[216] ; 
assign x0x2x3x5x6_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x5_share1 & x6_share1 ) ^ rand_bit[217] ; 
assign x0x2x3x5x6_subscript0_share2_1 = rand_bit[217] ; 
assign x1x2x3x4x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x4_share1 & x7_share1 ) ^ rand_bit[218] ; 
assign x1x2x3x4x7_subscript0_share2_1 = rand_bit[218] ; 
assign x0x1x2x3x4x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x4_share1 & x6_share1 ) ^ rand_bit[219] ; 
assign x0x1x2x3x4x6_subscript0_share2_1 = rand_bit[219] ; 
assign x0x1x2x3x4x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x4_share1 & x7_share1 ) ^ rand_bit[220] ; 
assign x0x1x2x3x4x7_subscript0_share2_1 = rand_bit[220] ; 
assign x0x1x2x3x5x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x5_share1 & x7_share1 ) ^ rand_bit[221] ; 
assign x0x1x2x3x5x7_subscript0_share2_1 = rand_bit[221] ; 
assign x0x1x2x3x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x6_share1 & x7_share1 ) ^ rand_bit[222] ; 
assign x0x1x2x3x6x7_subscript0_share2_1 = rand_bit[222] ; 
assign x0x1x2x4x5x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[223] ; 
assign x0x1x2x4x5x7_subscript0_share2_1 = rand_bit[223] ; 
assign x0x1x2x5x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[224] ; 
assign x0x1x2x5x6x7_subscript0_share2_1 = rand_bit[224] ; 
assign x0x1x3x4x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[225] ; 
assign x0x1x3x4x6x7_subscript0_share2_1 = rand_bit[225] ; 
assign x0x1x4x5x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[226] ; 
assign x0x1x4x5x6x7_subscript0_share2_1 = rand_bit[226] ; 
assign x0x2x3x4x5x6_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[227] ; 
assign x0x2x3x4x5x6_subscript0_share2_1 = rand_bit[227] ; 
assign x0x2x3x4x5x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[228] ; 
assign x0x2x3x4x5x7_subscript0_share2_1 = rand_bit[228] ; 
assign x0x2x3x5x6x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[229] ; 
assign x0x2x3x5x6x7_subscript0_share2_1 = rand_bit[229] ; 
assign x1x2x3x4x6x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[230] ; 
assign x1x2x3x4x6x7_subscript0_share2_1 = rand_bit[230] ; 
assign x1x2x4x5x6x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[231] ; 
assign x1x2x4x5x6x7_subscript0_share2_1 = rand_bit[231] ; 
assign x1x3x4x5x6x7_subscript0_share1_1 = ( x1_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[232] ; 
assign x1x3x4x5x6x7_subscript0_share2_1 = rand_bit[232] ; 
assign x2x3x4x5x6x7_subscript0_share1_1 = ( x2_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[233] ; 
assign x2x3x4x5x6x7_subscript0_share2_1 = rand_bit[233] ; 
assign x0x1x2x3x5x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x5_share1 & x6_share1 ) ^ rand_bit[234] ; 
assign x0x1x2x3x5x6_subscript0_share2_1 = rand_bit[234] ; 
assign x0x1x2x4x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[235] ; 
assign x0x1x2x4x6x7_subscript0_share2_1 = rand_bit[235] ; 
assign x0x1x3x4x5x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[236] ; 
assign x0x1x3x4x5x6_subscript0_share2_1 = rand_bit[236] ; 
assign x0x2x3x4x6x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[237] ; 
assign x0x2x3x4x6x7_subscript0_share2_1 = rand_bit[237] ; 
assign x1x2x3x4x5x6_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[238] ; 
assign x1x2x3x4x5x6_subscript0_share2_1 = rand_bit[238] ; 
assign x1x2x3x5x6x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[239] ; 
assign x1x2x3x5x6x7_subscript0_share2_1 = rand_bit[239] ; 
assign x0x1x2x3x4x5_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 ) ^ rand_bit[240] ; 
assign x0x1x2x3x4x5_subscript0_share2_1 = rand_bit[240] ; 
assign x0x1x2x4x5x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[241] ; 
assign x0x1x2x4x5x6_subscript0_share2_1 = rand_bit[241] ; 
assign x0x1x3x4x5x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[242] ; 
assign x0x1x3x4x5x7_subscript0_share2_1 = rand_bit[242] ; 
assign x0x1x3x5x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[243] ; 
assign x0x1x3x5x6x7_subscript0_share2_1 = rand_bit[243] ; 
assign x0x2x4x5x6x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[244] ; 
assign x0x2x4x5x6x7_subscript0_share2_1 = rand_bit[244] ; 
assign x1x2x3x4x5x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[245] ; 
assign x1x2x3x4x5x7_subscript0_share2_1 = rand_bit[245] ; 
assign x0x3x4x5x6x7_subscript0_share1_1 = ( x0_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[246] ; 
assign x0x3x4x5x6x7_subscript0_share2_1 = rand_bit[246] ; 
assign x0x1x2x3x4x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x4_share1 & x6_share1 & x7_share1 ) ^ rand_bit[247] ; 
assign x0x1x2x3x4x6x7_subscript0_share2_1 = rand_bit[247] ; 
assign x0x1x2x4x5x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[248] ; 
assign x0x1x2x4x5x6x7_subscript0_share2_1 = rand_bit[248] ; 
assign x0x2x3x4x5x6x7_subscript0_share1_1 = ( x0_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[249] ; 
assign x0x2x3x4x5x6x7_subscript0_share2_1 = rand_bit[249] ; 
assign x0x1x2x3x5x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[250] ; 
assign x0x1x2x3x5x6x7_subscript0_share2_1 = rand_bit[250] ; 
assign x0x1x3x4x5x6x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[251] ; 
assign x0x1x3x4x5x6x7_subscript0_share2_1 = rand_bit[251] ; 
assign x1x2x3x4x5x6x7_subscript0_share1_1 = ( x1_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 & x7_share1 ) ^ rand_bit[252] ; 
assign x1x2x3x4x5x6x7_subscript0_share2_1 = rand_bit[252] ; 
assign x0x1x2x3x4x5x6_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 & x6_share1 ) ^ rand_bit[253] ; 
assign x0x1x2x3x4x5x6_subscript0_share2_1 = rand_bit[253] ; 
assign x0x1x2x3x4x5x7_subscript0_share1_1 = ( x0_share1 & x1_share1 & x2_share1 & x3_share1 & x4_share1 & x5_share1 & x7_share1 ) ^ rand_bit[254] ; 
assign x0x1x2x3x4x5x7_subscript0_share2_1 = rand_bit[254] ; 


endmodule
