`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 02/22/2025
// Design Name: AES S-Box Two-Cycle First-Order Masked
// Module Name: AES_sbox_twocycle_firstorder
// Description: Implements a two-cycle first-order masked AES S-Box based on HO_TSM1.
// Dependencies: HO_TSM1 (First and Second Modules), sum_of_second_module_outputs, cross_module_multiplication, domain_inner
// Revision: 0.01 - Initial version
//////////////////////////////////////////////////////////////////////////////////

module AES_sbox_twocycle_firstorder ( clk, rand_bit,
	sbox_input_share1, sbox_input_share2,
    output_sbox_share1, output_sbox_share2
);


input clk;
input [46:1] rand_bit;


input [7:0] sbox_input_share1, sbox_input_share2;
output [7:0] output_sbox_share1, output_sbox_share2;


wire x0_input_share1 = sbox_input_share1[0];
wire x1_input_share1 = sbox_input_share1[1];
wire x2_input_share1 = sbox_input_share1[2];
wire x3_input_share1 = sbox_input_share1[3];
wire x4_input_share1 = sbox_input_share1[4];
wire x5_input_share1 = sbox_input_share1[5];
wire x6_input_share1 = sbox_input_share1[6];
wire x7_input_share1 = sbox_input_share1[7];

wire x0_input_share2 = sbox_input_share2[0];
wire x1_input_share2 = sbox_input_share2[1];
wire x2_input_share2 = sbox_input_share2[2];
wire x3_input_share2 = sbox_input_share2[3];
wire x4_input_share2 = sbox_input_share2[4];
wire x5_input_share2 = sbox_input_share2[5];
wire x6_input_share2 = sbox_input_share2[6];
wire x7_input_share2 = sbox_input_share2[7];

wire output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 ,    output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 ;
wire output_x4_share1, output_x5_share1, output_x6_share1, output_x7_share1, output_x4x5_share1, output_x4x6_share1, output_x4x7_share1, output_x5x6_share1, output_x5x7_share1, output_x6x7_share1, output_x4x5x6_share1, output_x4x5x7_share1, output_x4x6x7_share1, output_x5x6x7_share1, output_x4x5x6x7_share1 ,    output_x4_share2, output_x5_share2, output_x6_share2, output_x7_share2, output_x4x5_share2, output_x4x6_share2, output_x4x7_share2, output_x5x6_share2, output_x5x7_share2, output_x6x7_share2, output_x4x5x6_share2, output_x4x5x7_share2, output_x4x6x7_share2, output_x5x6x7_share2, output_x4x5x6x7_share2 ;

HO_TSM1 first_module(clk, rand_bit[19:1],   x0_input_share1, x1_input_share1, x2_input_share1, x3_input_share1,  x0_input_share2, x1_input_share2, x2_input_share2, x3_input_share2,    
output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 ,    output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 );
HO_TSM1 secon_module(clk, rand_bit[38:20],  x4_input_share1, x5_input_share1, x6_input_share1, x7_input_share1,  x4_input_share2, x5_input_share2, x6_input_share2, x7_input_share2,    
output_x4_share1, output_x5_share1, output_x6_share1, output_x7_share1, output_x4x5_share1, output_x4x6_share1, output_x4x7_share1, output_x5x6_share1, output_x5x7_share1, output_x6x7_share1, output_x4x5x6_share1, output_x4x5x7_share1, output_x4x6x7_share1, output_x5x6x7_share1, output_x4x5x6x7_share1 ,    output_x4_share2, output_x5_share2, output_x6_share2, output_x7_share2, output_x4x5_share2, output_x4x6_share2, output_x4x7_share2, output_x5x6_share2, output_x5x7_share2, output_x6x7_share2, output_x4x5x6_share2, output_x4x5x7_share2, output_x4x6x7_share2, output_x5x6x7_share2, output_x4x5x6x7_share2 );

wire [8:1] rand_bit_second;
assign rand_bit_second = rand_bit[46:39];



wire output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1 ;

wire output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2 ;

sum_of_second_module_outputs instance_share1 (
    output_x4_share1 ,  output_x5_share1 ,  output_x6_share1 ,  output_x7_share1 ,  output_x4x5_share1 ,  output_x4x6_share1 ,  output_x4x7_share1 ,  output_x5x6_share1 ,  output_x5x7_share1 ,  output_x6x7_share1 ,  output_x4x5x6_share1 ,  output_x4x5x7_share1 ,  output_x4x6x7_share1 ,  output_x5x6x7_share1 ,  output_x4x5x6x7_share1,
output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1

);

sum_of_second_module_outputs instance_share2 (
    output_x4_share2 ,  output_x5_share2 ,  output_x6_share2 ,  output_x7_share2 ,  output_x4x5_share2 ,  output_x4x6_share2 ,  output_x4x7_share2 ,  output_x5x6_share2 ,  output_x5x7_share2 ,  output_x6x7_share2 ,  output_x4x5x6_share2 ,  output_x4x5x7_share2 ,  output_x4x6x7_share2 ,  output_x5x6x7_share2 ,  output_x4x5x6x7_share2,
output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2

);



wire cross_module_equation_num0_domain_1, cross_module_equation_num1_domain_1, cross_module_equation_num2_domain_1, cross_module_equation_num3_domain_1,cross_module_equation_num4_domain_1,cross_module_equation_num5_domain_1,cross_module_equation_num6_domain_1,cross_module_equation_num7_domain_1;
wire cross_module_equation_num0_domain_2, cross_module_equation_num1_domain_2, cross_module_equation_num2_domain_2, cross_module_equation_num3_domain_2,cross_module_equation_num4_domain_2,cross_module_equation_num5_domain_2,cross_module_equation_num6_domain_2,cross_module_equation_num7_domain_2;
wire cross_module_equation_num0_domain_3, cross_module_equation_num1_domain_3, cross_module_equation_num2_domain_3, cross_module_equation_num3_domain_3,cross_module_equation_num4_domain_3,cross_module_equation_num5_domain_3,cross_module_equation_num6_domain_3,cross_module_equation_num7_domain_3;
wire cross_module_equation_num0_domain_4, cross_module_equation_num1_domain_4, cross_module_equation_num2_domain_4, cross_module_equation_num3_domain_4,cross_module_equation_num4_domain_4,cross_module_equation_num5_domain_4,cross_module_equation_num6_domain_4,cross_module_equation_num7_domain_4;


cross_module_multiplication inst1 (
output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 , 
output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1,
cross_module_equation_num0_domain_1, cross_module_equation_num1_domain_1, cross_module_equation_num2_domain_1, cross_module_equation_num3_domain_1,cross_module_equation_num4_domain_1,cross_module_equation_num5_domain_1,cross_module_equation_num6_domain_1,cross_module_equation_num7_domain_1
);


cross_module_multiplication inst2 (
output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 , 
output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2,
cross_module_equation_num0_domain_2, cross_module_equation_num1_domain_2, cross_module_equation_num2_domain_2, cross_module_equation_num3_domain_2,cross_module_equation_num4_domain_2,cross_module_equation_num5_domain_2,cross_module_equation_num6_domain_2,cross_module_equation_num7_domain_2
);

cross_module_multiplication inst3 (
output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 , 
output_sum_secondmodule_equation_num_0_index_0_share1, output_sum_secondmodule_equation_num_0_index_1_share1, output_sum_secondmodule_equation_num_0_index_2_share1, output_sum_secondmodule_equation_num_0_index_3_share1, output_sum_secondmodule_equation_num_0_index_4_share1, output_sum_secondmodule_equation_num_0_index_5_share1, output_sum_secondmodule_equation_num_0_index_6_share1, output_sum_secondmodule_equation_num_0_index_7_share1, output_sum_secondmodule_equation_num_0_index_8_share1, output_sum_secondmodule_equation_num_0_index_9_share1, output_sum_secondmodule_equation_num_0_index_10_share1, output_sum_secondmodule_equation_num_0_index_11_share1, output_sum_secondmodule_equation_num_0_index_12_share1, output_sum_secondmodule_equation_num_0_index_13_share1, output_sum_secondmodule_equation_num_0_index_14_share1,
output_sum_secondmodule_equation_num_1_index_0_share1, output_sum_secondmodule_equation_num_1_index_1_share1, output_sum_secondmodule_equation_num_1_index_2_share1, output_sum_secondmodule_equation_num_1_index_3_share1, output_sum_secondmodule_equation_num_1_index_4_share1, output_sum_secondmodule_equation_num_1_index_5_share1, output_sum_secondmodule_equation_num_1_index_6_share1, output_sum_secondmodule_equation_num_1_index_7_share1, output_sum_secondmodule_equation_num_1_index_8_share1, output_sum_secondmodule_equation_num_1_index_9_share1, output_sum_secondmodule_equation_num_1_index_10_share1, output_sum_secondmodule_equation_num_1_index_11_share1, output_sum_secondmodule_equation_num_1_index_12_share1, output_sum_secondmodule_equation_num_1_index_13_share1, output_sum_secondmodule_equation_num_1_index_14_share1,
output_sum_secondmodule_equation_num_2_index_0_share1, output_sum_secondmodule_equation_num_2_index_1_share1, output_sum_secondmodule_equation_num_2_index_2_share1, output_sum_secondmodule_equation_num_2_index_3_share1, output_sum_secondmodule_equation_num_2_index_4_share1, output_sum_secondmodule_equation_num_2_index_5_share1, output_sum_secondmodule_equation_num_2_index_6_share1, output_sum_secondmodule_equation_num_2_index_7_share1, output_sum_secondmodule_equation_num_2_index_8_share1, output_sum_secondmodule_equation_num_2_index_9_share1, output_sum_secondmodule_equation_num_2_index_10_share1, output_sum_secondmodule_equation_num_2_index_11_share1, output_sum_secondmodule_equation_num_2_index_12_share1, output_sum_secondmodule_equation_num_2_index_13_share1, output_sum_secondmodule_equation_num_2_index_14_share1,
output_sum_secondmodule_equation_num_3_index_0_share1, output_sum_secondmodule_equation_num_3_index_1_share1, output_sum_secondmodule_equation_num_3_index_2_share1, output_sum_secondmodule_equation_num_3_index_3_share1, output_sum_secondmodule_equation_num_3_index_4_share1, output_sum_secondmodule_equation_num_3_index_5_share1, output_sum_secondmodule_equation_num_3_index_6_share1, output_sum_secondmodule_equation_num_3_index_7_share1, output_sum_secondmodule_equation_num_3_index_8_share1, output_sum_secondmodule_equation_num_3_index_9_share1, output_sum_secondmodule_equation_num_3_index_10_share1, output_sum_secondmodule_equation_num_3_index_11_share1, output_sum_secondmodule_equation_num_3_index_12_share1, output_sum_secondmodule_equation_num_3_index_13_share1, output_sum_secondmodule_equation_num_3_index_14_share1,
output_sum_secondmodule_equation_num_4_index_0_share1, output_sum_secondmodule_equation_num_4_index_1_share1, output_sum_secondmodule_equation_num_4_index_2_share1, output_sum_secondmodule_equation_num_4_index_3_share1, output_sum_secondmodule_equation_num_4_index_4_share1, output_sum_secondmodule_equation_num_4_index_5_share1, output_sum_secondmodule_equation_num_4_index_6_share1, output_sum_secondmodule_equation_num_4_index_7_share1, output_sum_secondmodule_equation_num_4_index_8_share1, output_sum_secondmodule_equation_num_4_index_9_share1, output_sum_secondmodule_equation_num_4_index_10_share1, output_sum_secondmodule_equation_num_4_index_11_share1, output_sum_secondmodule_equation_num_4_index_12_share1, output_sum_secondmodule_equation_num_4_index_13_share1, output_sum_secondmodule_equation_num_4_index_14_share1,
output_sum_secondmodule_equation_num_5_index_0_share1, output_sum_secondmodule_equation_num_5_index_1_share1, output_sum_secondmodule_equation_num_5_index_2_share1, output_sum_secondmodule_equation_num_5_index_3_share1, output_sum_secondmodule_equation_num_5_index_4_share1, output_sum_secondmodule_equation_num_5_index_5_share1, output_sum_secondmodule_equation_num_5_index_6_share1, output_sum_secondmodule_equation_num_5_index_7_share1, output_sum_secondmodule_equation_num_5_index_8_share1, output_sum_secondmodule_equation_num_5_index_9_share1, output_sum_secondmodule_equation_num_5_index_10_share1, output_sum_secondmodule_equation_num_5_index_11_share1, output_sum_secondmodule_equation_num_5_index_12_share1, output_sum_secondmodule_equation_num_5_index_13_share1, output_sum_secondmodule_equation_num_5_index_14_share1,
output_sum_secondmodule_equation_num_6_index_0_share1, output_sum_secondmodule_equation_num_6_index_1_share1, output_sum_secondmodule_equation_num_6_index_2_share1, output_sum_secondmodule_equation_num_6_index_3_share1, output_sum_secondmodule_equation_num_6_index_4_share1, output_sum_secondmodule_equation_num_6_index_5_share1, output_sum_secondmodule_equation_num_6_index_6_share1, output_sum_secondmodule_equation_num_6_index_7_share1, output_sum_secondmodule_equation_num_6_index_8_share1, output_sum_secondmodule_equation_num_6_index_9_share1, output_sum_secondmodule_equation_num_6_index_10_share1, output_sum_secondmodule_equation_num_6_index_11_share1, output_sum_secondmodule_equation_num_6_index_12_share1, output_sum_secondmodule_equation_num_6_index_13_share1, output_sum_secondmodule_equation_num_6_index_14_share1,
output_sum_secondmodule_equation_num_7_index_0_share1, output_sum_secondmodule_equation_num_7_index_1_share1, output_sum_secondmodule_equation_num_7_index_2_share1, output_sum_secondmodule_equation_num_7_index_3_share1, output_sum_secondmodule_equation_num_7_index_4_share1, output_sum_secondmodule_equation_num_7_index_5_share1, output_sum_secondmodule_equation_num_7_index_6_share1, output_sum_secondmodule_equation_num_7_index_7_share1, output_sum_secondmodule_equation_num_7_index_8_share1, output_sum_secondmodule_equation_num_7_index_9_share1, output_sum_secondmodule_equation_num_7_index_10_share1, output_sum_secondmodule_equation_num_7_index_11_share1, output_sum_secondmodule_equation_num_7_index_12_share1, output_sum_secondmodule_equation_num_7_index_13_share1, output_sum_secondmodule_equation_num_7_index_14_share1,
cross_module_equation_num0_domain_3, cross_module_equation_num1_domain_3, cross_module_equation_num2_domain_3, cross_module_equation_num3_domain_3,cross_module_equation_num4_domain_3,cross_module_equation_num5_domain_3,cross_module_equation_num6_domain_3,cross_module_equation_num7_domain_3
);

cross_module_multiplication inst4 (
output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 , 
output_sum_secondmodule_equation_num_0_index_0_share2, output_sum_secondmodule_equation_num_0_index_1_share2, output_sum_secondmodule_equation_num_0_index_2_share2, output_sum_secondmodule_equation_num_0_index_3_share2, output_sum_secondmodule_equation_num_0_index_4_share2, output_sum_secondmodule_equation_num_0_index_5_share2, output_sum_secondmodule_equation_num_0_index_6_share2, output_sum_secondmodule_equation_num_0_index_7_share2, output_sum_secondmodule_equation_num_0_index_8_share2, output_sum_secondmodule_equation_num_0_index_9_share2, output_sum_secondmodule_equation_num_0_index_10_share2, output_sum_secondmodule_equation_num_0_index_11_share2, output_sum_secondmodule_equation_num_0_index_12_share2, output_sum_secondmodule_equation_num_0_index_13_share2, output_sum_secondmodule_equation_num_0_index_14_share2,
output_sum_secondmodule_equation_num_1_index_0_share2, output_sum_secondmodule_equation_num_1_index_1_share2, output_sum_secondmodule_equation_num_1_index_2_share2, output_sum_secondmodule_equation_num_1_index_3_share2, output_sum_secondmodule_equation_num_1_index_4_share2, output_sum_secondmodule_equation_num_1_index_5_share2, output_sum_secondmodule_equation_num_1_index_6_share2, output_sum_secondmodule_equation_num_1_index_7_share2, output_sum_secondmodule_equation_num_1_index_8_share2, output_sum_secondmodule_equation_num_1_index_9_share2, output_sum_secondmodule_equation_num_1_index_10_share2, output_sum_secondmodule_equation_num_1_index_11_share2, output_sum_secondmodule_equation_num_1_index_12_share2, output_sum_secondmodule_equation_num_1_index_13_share2, output_sum_secondmodule_equation_num_1_index_14_share2,
output_sum_secondmodule_equation_num_2_index_0_share2, output_sum_secondmodule_equation_num_2_index_1_share2, output_sum_secondmodule_equation_num_2_index_2_share2, output_sum_secondmodule_equation_num_2_index_3_share2, output_sum_secondmodule_equation_num_2_index_4_share2, output_sum_secondmodule_equation_num_2_index_5_share2, output_sum_secondmodule_equation_num_2_index_6_share2, output_sum_secondmodule_equation_num_2_index_7_share2, output_sum_secondmodule_equation_num_2_index_8_share2, output_sum_secondmodule_equation_num_2_index_9_share2, output_sum_secondmodule_equation_num_2_index_10_share2, output_sum_secondmodule_equation_num_2_index_11_share2, output_sum_secondmodule_equation_num_2_index_12_share2, output_sum_secondmodule_equation_num_2_index_13_share2, output_sum_secondmodule_equation_num_2_index_14_share2,
output_sum_secondmodule_equation_num_3_index_0_share2, output_sum_secondmodule_equation_num_3_index_1_share2, output_sum_secondmodule_equation_num_3_index_2_share2, output_sum_secondmodule_equation_num_3_index_3_share2, output_sum_secondmodule_equation_num_3_index_4_share2, output_sum_secondmodule_equation_num_3_index_5_share2, output_sum_secondmodule_equation_num_3_index_6_share2, output_sum_secondmodule_equation_num_3_index_7_share2, output_sum_secondmodule_equation_num_3_index_8_share2, output_sum_secondmodule_equation_num_3_index_9_share2, output_sum_secondmodule_equation_num_3_index_10_share2, output_sum_secondmodule_equation_num_3_index_11_share2, output_sum_secondmodule_equation_num_3_index_12_share2, output_sum_secondmodule_equation_num_3_index_13_share2, output_sum_secondmodule_equation_num_3_index_14_share2,
output_sum_secondmodule_equation_num_4_index_0_share2, output_sum_secondmodule_equation_num_4_index_1_share2, output_sum_secondmodule_equation_num_4_index_2_share2, output_sum_secondmodule_equation_num_4_index_3_share2, output_sum_secondmodule_equation_num_4_index_4_share2, output_sum_secondmodule_equation_num_4_index_5_share2, output_sum_secondmodule_equation_num_4_index_6_share2, output_sum_secondmodule_equation_num_4_index_7_share2, output_sum_secondmodule_equation_num_4_index_8_share2, output_sum_secondmodule_equation_num_4_index_9_share2, output_sum_secondmodule_equation_num_4_index_10_share2, output_sum_secondmodule_equation_num_4_index_11_share2, output_sum_secondmodule_equation_num_4_index_12_share2, output_sum_secondmodule_equation_num_4_index_13_share2, output_sum_secondmodule_equation_num_4_index_14_share2,
output_sum_secondmodule_equation_num_5_index_0_share2, output_sum_secondmodule_equation_num_5_index_1_share2, output_sum_secondmodule_equation_num_5_index_2_share2, output_sum_secondmodule_equation_num_5_index_3_share2, output_sum_secondmodule_equation_num_5_index_4_share2, output_sum_secondmodule_equation_num_5_index_5_share2, output_sum_secondmodule_equation_num_5_index_6_share2, output_sum_secondmodule_equation_num_5_index_7_share2, output_sum_secondmodule_equation_num_5_index_8_share2, output_sum_secondmodule_equation_num_5_index_9_share2, output_sum_secondmodule_equation_num_5_index_10_share2, output_sum_secondmodule_equation_num_5_index_11_share2, output_sum_secondmodule_equation_num_5_index_12_share2, output_sum_secondmodule_equation_num_5_index_13_share2, output_sum_secondmodule_equation_num_5_index_14_share2,
output_sum_secondmodule_equation_num_6_index_0_share2, output_sum_secondmodule_equation_num_6_index_1_share2, output_sum_secondmodule_equation_num_6_index_2_share2, output_sum_secondmodule_equation_num_6_index_3_share2, output_sum_secondmodule_equation_num_6_index_4_share2, output_sum_secondmodule_equation_num_6_index_5_share2, output_sum_secondmodule_equation_num_6_index_6_share2, output_sum_secondmodule_equation_num_6_index_7_share2, output_sum_secondmodule_equation_num_6_index_8_share2, output_sum_secondmodule_equation_num_6_index_9_share2, output_sum_secondmodule_equation_num_6_index_10_share2, output_sum_secondmodule_equation_num_6_index_11_share2, output_sum_secondmodule_equation_num_6_index_12_share2, output_sum_secondmodule_equation_num_6_index_13_share2, output_sum_secondmodule_equation_num_6_index_14_share2,
output_sum_secondmodule_equation_num_7_index_0_share2, output_sum_secondmodule_equation_num_7_index_1_share2, output_sum_secondmodule_equation_num_7_index_2_share2, output_sum_secondmodule_equation_num_7_index_3_share2, output_sum_secondmodule_equation_num_7_index_4_share2, output_sum_secondmodule_equation_num_7_index_5_share2, output_sum_secondmodule_equation_num_7_index_6_share2, output_sum_secondmodule_equation_num_7_index_7_share2, output_sum_secondmodule_equation_num_7_index_8_share2, output_sum_secondmodule_equation_num_7_index_9_share2, output_sum_secondmodule_equation_num_7_index_10_share2, output_sum_secondmodule_equation_num_7_index_11_share2, output_sum_secondmodule_equation_num_7_index_12_share2, output_sum_secondmodule_equation_num_7_index_13_share2, output_sum_secondmodule_equation_num_7_index_14_share2,
cross_module_equation_num0_domain_4, cross_module_equation_num1_domain_4, cross_module_equation_num2_domain_4, cross_module_equation_num3_domain_4,cross_module_equation_num4_domain_4,cross_module_equation_num5_domain_4,cross_module_equation_num6_domain_4,cross_module_equation_num7_domain_4
);

wire inner_module_equation_num0_domain_1 , inner_module_equation_num1_domain_1 , inner_module_equation_num2_domain_1 , inner_module_equation_num3_domain_1 , inner_module_equation_num4_domain_1 , inner_module_equation_num5_domain_1 , inner_module_equation_num6_domain_1 , inner_module_equation_num7_domain_1 ;
wire inner_module_equation_num0_domain_4 , inner_module_equation_num1_domain_4 , inner_module_equation_num2_domain_4 , inner_module_equation_num3_domain_4 , inner_module_equation_num4_domain_4 , inner_module_equation_num5_domain_4 , inner_module_equation_num6_domain_4 , inner_module_equation_num7_domain_4 ;

domain_inner domain1_inst(   output_x0_share1, output_x1_share1, output_x2_share1, output_x3_share1, output_x0x1_share1, output_x0x2_share1, output_x0x3_share1, output_x1x2_share1, output_x1x3_share1, output_x2x3_share1, output_x0x1x2_share1, output_x0x1x3_share1, output_x0x2x3_share1, output_x1x2x3_share1, output_x0x1x2x3_share1 ,   output_x4_share1, output_x5_share1, output_x6_share1, output_x7_share1, output_x4x5_share1, output_x4x6_share1, output_x4x7_share1, output_x5x6_share1, output_x5x7_share1, output_x6x7_share1, output_x4x5x6_share1, output_x4x5x7_share1, output_x4x6x7_share1, output_x5x6x7_share1, output_x4x5x6x7_share1 , 
inner_module_equation_num0_domain_1 , inner_module_equation_num1_domain_1 , inner_module_equation_num2_domain_1 , inner_module_equation_num3_domain_1 , inner_module_equation_num4_domain_1 , inner_module_equation_num5_domain_1 , inner_module_equation_num6_domain_1 , inner_module_equation_num7_domain_1 );

domain_inner domain4_inst(   output_x0_share2, output_x1_share2, output_x2_share2, output_x3_share2, output_x0x1_share2, output_x0x2_share2, output_x0x3_share2, output_x1x2_share2, output_x1x3_share2, output_x2x3_share2, output_x0x1x2_share2, output_x0x1x3_share2, output_x0x2x3_share2, output_x1x2x3_share2, output_x0x1x2x3_share2 ,   output_x4_share2, output_x5_share2, output_x6_share2, output_x7_share2, output_x4x5_share2, output_x4x6_share2, output_x4x7_share2, output_x5x6_share2, output_x5x7_share2, output_x6x7_share2, output_x4x5x6_share2, output_x4x5x7_share2, output_x4x6x7_share2, output_x5x6x7_share2, output_x4x5x6x7_share2 , 
inner_module_equation_num0_domain_4 , inner_module_equation_num1_domain_4 , inner_module_equation_num2_domain_4 , inner_module_equation_num3_domain_4 , inner_module_equation_num4_domain_4 , inner_module_equation_num5_domain_4 , inner_module_equation_num6_domain_4 , inner_module_equation_num7_domain_4 );

wire inner_module_equation_num0_domain_2 ;
wire inner_module_equation_num1_domain_2 ;
wire inner_module_equation_num2_domain_2 ;
wire inner_module_equation_num3_domain_2 ;
wire inner_module_equation_num4_domain_2 ;
wire inner_module_equation_num5_domain_2 ;
wire inner_module_equation_num6_domain_2 ;
wire inner_module_equation_num7_domain_2 ;

assign inner_module_equation_num0_domain_2= 1'b0 ;
assign inner_module_equation_num1_domain_2= 1'b0 ;
assign inner_module_equation_num2_domain_2= 1'b0 ;
assign inner_module_equation_num3_domain_2= 1'b0 ;
assign inner_module_equation_num4_domain_2= 1'b0 ;
assign inner_module_equation_num5_domain_2= 1'b0 ;
assign inner_module_equation_num6_domain_2= 1'b0 ;
assign inner_module_equation_num7_domain_2= 1'b0 ;

wire inner_module_equation_num0_domain_3 ;
wire inner_module_equation_num1_domain_3 ;
wire inner_module_equation_num2_domain_3 ;
wire inner_module_equation_num3_domain_3 ;
wire inner_module_equation_num4_domain_3 ;
wire inner_module_equation_num5_domain_3 ;
wire inner_module_equation_num6_domain_3 ;
wire inner_module_equation_num7_domain_3 ;

assign inner_module_equation_num0_domain_3= 1'b0 ;
assign inner_module_equation_num1_domain_3= 1'b0 ;
assign inner_module_equation_num2_domain_3= 1'b0 ;
assign inner_module_equation_num3_domain_3= 1'b0 ;
assign inner_module_equation_num4_domain_3= 1'b0 ;
assign inner_module_equation_num5_domain_3= 1'b0 ;
assign inner_module_equation_num6_domain_3= 1'b0 ;
assign inner_module_equation_num7_domain_3= 1'b0 ;

wire inner_plus_cross_module_equation_num0_domain_1, inner_plus_cross_module_equation_num0_domain_2, inner_plus_cross_module_equation_num0_domain_3, inner_plus_cross_module_equation_num0_domain_4;
wire inner_plus_cross_module_equation_num1_domain_1, inner_plus_cross_module_equation_num1_domain_2, inner_plus_cross_module_equation_num1_domain_3, inner_plus_cross_module_equation_num1_domain_4;
wire inner_plus_cross_module_equation_num2_domain_1, inner_plus_cross_module_equation_num2_domain_2, inner_plus_cross_module_equation_num2_domain_3, inner_plus_cross_module_equation_num2_domain_4;
wire inner_plus_cross_module_equation_num3_domain_1, inner_plus_cross_module_equation_num3_domain_2, inner_plus_cross_module_equation_num3_domain_3, inner_plus_cross_module_equation_num3_domain_4;
wire inner_plus_cross_module_equation_num4_domain_1, inner_plus_cross_module_equation_num4_domain_2, inner_plus_cross_module_equation_num4_domain_3, inner_plus_cross_module_equation_num4_domain_4;
wire inner_plus_cross_module_equation_num5_domain_1, inner_plus_cross_module_equation_num5_domain_2, inner_plus_cross_module_equation_num5_domain_3, inner_plus_cross_module_equation_num5_domain_4;
wire inner_plus_cross_module_equation_num6_domain_1, inner_plus_cross_module_equation_num6_domain_2, inner_plus_cross_module_equation_num6_domain_3, inner_plus_cross_module_equation_num6_domain_4;
wire inner_plus_cross_module_equation_num7_domain_1, inner_plus_cross_module_equation_num7_domain_2, inner_plus_cross_module_equation_num7_domain_3, inner_plus_cross_module_equation_num7_domain_4;


xor_module xor_num0_dom1(cross_module_equation_num0_domain_1,inner_module_equation_num0_domain_1,inner_plus_cross_module_equation_num0_domain_1);
xor_module xor_num0_dom2(cross_module_equation_num0_domain_2,inner_module_equation_num0_domain_2,inner_plus_cross_module_equation_num0_domain_2);
xor_module xor_num0_dom3(cross_module_equation_num0_domain_3,inner_module_equation_num0_domain_3,inner_plus_cross_module_equation_num0_domain_3);
xor_module xor_num0_dom4(cross_module_equation_num0_domain_4,inner_module_equation_num0_domain_4,inner_plus_cross_module_equation_num0_domain_4);

xor_module xor_num1_dom1(cross_module_equation_num1_domain_1,inner_module_equation_num1_domain_1,inner_plus_cross_module_equation_num1_domain_1);
xor_module xor_num1_dom2(cross_module_equation_num1_domain_2,inner_module_equation_num1_domain_2,inner_plus_cross_module_equation_num1_domain_2);
xor_module xor_num1_dom3(cross_module_equation_num1_domain_3,inner_module_equation_num1_domain_3,inner_plus_cross_module_equation_num1_domain_3);
xor_module xor_num1_dom4(cross_module_equation_num1_domain_4,inner_module_equation_num1_domain_4,inner_plus_cross_module_equation_num1_domain_4);

xor_module xor_num2_dom1(cross_module_equation_num2_domain_1,inner_module_equation_num2_domain_1,inner_plus_cross_module_equation_num2_domain_1);
xor_module xor_num2_dom2(cross_module_equation_num2_domain_2,inner_module_equation_num2_domain_2,inner_plus_cross_module_equation_num2_domain_2);
xor_module xor_num2_dom3(cross_module_equation_num2_domain_3,inner_module_equation_num2_domain_3,inner_plus_cross_module_equation_num2_domain_3);
xor_module xor_num2_dom4(cross_module_equation_num2_domain_4,inner_module_equation_num2_domain_4,inner_plus_cross_module_equation_num2_domain_4);

xor_module xor_num3_dom1(cross_module_equation_num3_domain_1,inner_module_equation_num3_domain_1,inner_plus_cross_module_equation_num3_domain_1);
xor_module xor_num3_dom2(cross_module_equation_num3_domain_2,inner_module_equation_num3_domain_2,inner_plus_cross_module_equation_num3_domain_2);
xor_module xor_num3_dom3(cross_module_equation_num3_domain_3,inner_module_equation_num3_domain_3,inner_plus_cross_module_equation_num3_domain_3);
xor_module xor_num3_dom4(cross_module_equation_num3_domain_4,inner_module_equation_num3_domain_4,inner_plus_cross_module_equation_num3_domain_4);

xor_module xor_num4_dom1(cross_module_equation_num4_domain_1,inner_module_equation_num4_domain_1,inner_plus_cross_module_equation_num4_domain_1);
xor_module xor_num4_dom2(cross_module_equation_num4_domain_2,inner_module_equation_num4_domain_2,inner_plus_cross_module_equation_num4_domain_2);
xor_module xor_num4_dom3(cross_module_equation_num4_domain_3,inner_module_equation_num4_domain_3,inner_plus_cross_module_equation_num4_domain_3);
xor_module xor_num4_dom4(cross_module_equation_num4_domain_4,inner_module_equation_num4_domain_4,inner_plus_cross_module_equation_num4_domain_4);

xor_module xor_num5_dom1(cross_module_equation_num5_domain_1,inner_module_equation_num5_domain_1,inner_plus_cross_module_equation_num5_domain_1);
xor_module xor_num5_dom2(cross_module_equation_num5_domain_2,inner_module_equation_num5_domain_2,inner_plus_cross_module_equation_num5_domain_2);
xor_module xor_num5_dom3(cross_module_equation_num5_domain_3,inner_module_equation_num5_domain_3,inner_plus_cross_module_equation_num5_domain_3);
xor_module xor_num5_dom4(cross_module_equation_num5_domain_4,inner_module_equation_num5_domain_4,inner_plus_cross_module_equation_num5_domain_4);

xor_module xor_num6_dom1(cross_module_equation_num6_domain_1,inner_module_equation_num6_domain_1,inner_plus_cross_module_equation_num6_domain_1);
xor_module xor_num6_dom2(cross_module_equation_num6_domain_2,inner_module_equation_num6_domain_2,inner_plus_cross_module_equation_num6_domain_2);
xor_module xor_num6_dom3(cross_module_equation_num6_domain_3,inner_module_equation_num6_domain_3,inner_plus_cross_module_equation_num6_domain_3);
xor_module xor_num6_dom4(cross_module_equation_num6_domain_4,inner_module_equation_num6_domain_4,inner_plus_cross_module_equation_num6_domain_4);

xor_module xor_num7_dom1(cross_module_equation_num7_domain_1,inner_module_equation_num7_domain_1,inner_plus_cross_module_equation_num7_domain_1);
xor_module xor_num7_dom2(cross_module_equation_num7_domain_2,inner_module_equation_num7_domain_2,inner_plus_cross_module_equation_num7_domain_2);
xor_module xor_num7_dom3(cross_module_equation_num7_domain_3,inner_module_equation_num7_domain_3,inner_plus_cross_module_equation_num7_domain_3);
xor_module xor_num7_dom4(cross_module_equation_num7_domain_4,inner_module_equation_num7_domain_4,inner_plus_cross_module_equation_num7_domain_4);





reg sbox_out_num_0_domain_1_reg,sbox_out_num_0_domain_2_reg,sbox_out_num_0_domain_3_reg,sbox_out_num_0_domain_4_reg ;
always@(posedge clk)
begin
	sbox_out_num_0_domain_1_reg <= inner_plus_cross_module_equation_num0_domain_1 ^ 1'b1;
	sbox_out_num_0_domain_2_reg <= inner_plus_cross_module_equation_num0_domain_2 ^ rand_bit_second[1] ;
	sbox_out_num_0_domain_3_reg <= inner_plus_cross_module_equation_num0_domain_3 ^ rand_bit_second[1] ;
	sbox_out_num_0_domain_4_reg <= inner_plus_cross_module_equation_num0_domain_4 ;
end

wire sbox_out_num_0_share1, sbox_out_num_0_share2 ;
assign sbox_out_num_0_share1 = sbox_out_num_0_domain_1_reg ^ sbox_out_num_0_domain_2_reg ;
assign sbox_out_num_0_share2 = sbox_out_num_0_domain_3_reg ^ sbox_out_num_0_domain_4_reg ;



reg sbox_out_num_1_domain_1_reg,sbox_out_num_1_domain_2_reg,sbox_out_num_1_domain_3_reg,sbox_out_num_1_domain_4_reg ;
always@(posedge clk)
begin
	sbox_out_num_1_domain_1_reg <= inner_plus_cross_module_equation_num1_domain_1 ^ 1'b1;
	sbox_out_num_1_domain_2_reg <= inner_plus_cross_module_equation_num1_domain_2 ^ rand_bit_second[2] ;
	sbox_out_num_1_domain_3_reg <= inner_plus_cross_module_equation_num1_domain_3 ^ rand_bit_second[2] ;
	sbox_out_num_1_domain_4_reg <= inner_plus_cross_module_equation_num1_domain_4 ;
end

wire sbox_out_num_1_share1, sbox_out_num_1_share2 ;
assign sbox_out_num_1_share1 = sbox_out_num_1_domain_1_reg ^ sbox_out_num_1_domain_2_reg ;
assign sbox_out_num_1_share2 = sbox_out_num_1_domain_3_reg ^ sbox_out_num_1_domain_4_reg ;



reg sbox_out_num_2_domain_1_reg,sbox_out_num_2_domain_2_reg,sbox_out_num_2_domain_3_reg,sbox_out_num_2_domain_4_reg ;
always@(posedge clk)
begin
	sbox_out_num_2_domain_1_reg <= inner_plus_cross_module_equation_num2_domain_1 ;
	sbox_out_num_2_domain_2_reg <= inner_plus_cross_module_equation_num2_domain_2 ^ rand_bit_second[3] ;
	sbox_out_num_2_domain_3_reg <= inner_plus_cross_module_equation_num2_domain_3 ^ rand_bit_second[3] ;
	sbox_out_num_2_domain_4_reg <= inner_plus_cross_module_equation_num2_domain_4 ;
end

wire sbox_out_num_2_share1, sbox_out_num_2_share2 ;
assign sbox_out_num_2_share1 = sbox_out_num_2_domain_1_reg ^ sbox_out_num_2_domain_2_reg ;
assign sbox_out_num_2_share2 = sbox_out_num_2_domain_3_reg ^ sbox_out_num_2_domain_4_reg ;



reg sbox_out_num_3_domain_1_reg,sbox_out_num_3_domain_2_reg,sbox_out_num_3_domain_3_reg,sbox_out_num_3_domain_4_reg ;
always@(posedge clk)
begin
	sbox_out_num_3_domain_1_reg <= inner_plus_cross_module_equation_num3_domain_1 ;
	sbox_out_num_3_domain_2_reg <= inner_plus_cross_module_equation_num3_domain_2 ^ rand_bit_second[4] ;
	sbox_out_num_3_domain_3_reg <= inner_plus_cross_module_equation_num3_domain_3 ^ rand_bit_second[4] ;
	sbox_out_num_3_domain_4_reg <= inner_plus_cross_module_equation_num3_domain_4 ;
end

wire sbox_out_num_3_share1, sbox_out_num_3_share2 ;
assign sbox_out_num_3_share1 = sbox_out_num_3_domain_1_reg ^ sbox_out_num_3_domain_2_reg ;
assign sbox_out_num_3_share2 = sbox_out_num_3_domain_3_reg ^ sbox_out_num_3_domain_4_reg ;



reg sbox_out_num_4_domain_1_reg,sbox_out_num_4_domain_2_reg,sbox_out_num_4_domain_3_reg,sbox_out_num_4_domain_4_reg ;
always@(posedge clk)
begin
	sbox_out_num_4_domain_1_reg <= inner_plus_cross_module_equation_num4_domain_1 ;
	sbox_out_num_4_domain_2_reg <= inner_plus_cross_module_equation_num4_domain_2 ^ rand_bit_second[5] ;
	sbox_out_num_4_domain_3_reg <= inner_plus_cross_module_equation_num4_domain_3 ^ rand_bit_second[5] ;
	sbox_out_num_4_domain_4_reg <= inner_plus_cross_module_equation_num4_domain_4 ;
end

wire sbox_out_num_4_share1, sbox_out_num_4_share2 ;
assign sbox_out_num_4_share1 = sbox_out_num_4_domain_1_reg ^ sbox_out_num_4_domain_2_reg ;
assign sbox_out_num_4_share2 = sbox_out_num_4_domain_3_reg ^ sbox_out_num_4_domain_4_reg ;



reg sbox_out_num_5_domain_1_reg,sbox_out_num_5_domain_2_reg,sbox_out_num_5_domain_3_reg,sbox_out_num_5_domain_4_reg ;
always@(posedge clk)
begin
	sbox_out_num_5_domain_1_reg <= inner_plus_cross_module_equation_num5_domain_1 ^ 1'b1;
	sbox_out_num_5_domain_2_reg <= inner_plus_cross_module_equation_num5_domain_2 ^ rand_bit_second[6] ;
	sbox_out_num_5_domain_3_reg <= inner_plus_cross_module_equation_num5_domain_3 ^ rand_bit_second[6] ;
	sbox_out_num_5_domain_4_reg <= inner_plus_cross_module_equation_num5_domain_4 ;
end

wire sbox_out_num_5_share1, sbox_out_num_5_share2 ;
assign sbox_out_num_5_share1 = sbox_out_num_5_domain_1_reg ^ sbox_out_num_5_domain_2_reg ;
assign sbox_out_num_5_share2 = sbox_out_num_5_domain_3_reg ^ sbox_out_num_5_domain_4_reg ;



reg sbox_out_num_6_domain_1_reg,sbox_out_num_6_domain_2_reg,sbox_out_num_6_domain_3_reg,sbox_out_num_6_domain_4_reg ;
always@(posedge clk)
begin
	sbox_out_num_6_domain_1_reg <= inner_plus_cross_module_equation_num6_domain_1 ^ 1'b1;
	sbox_out_num_6_domain_2_reg <= inner_plus_cross_module_equation_num6_domain_2 ^ rand_bit_second[7] ;
	sbox_out_num_6_domain_3_reg <= inner_plus_cross_module_equation_num6_domain_3 ^ rand_bit_second[7] ;
	sbox_out_num_6_domain_4_reg <= inner_plus_cross_module_equation_num6_domain_4 ;
end

wire sbox_out_num_6_share1, sbox_out_num_6_share2 ;
assign sbox_out_num_6_share1 = sbox_out_num_6_domain_1_reg ^ sbox_out_num_6_domain_2_reg ;
assign sbox_out_num_6_share2 = sbox_out_num_6_domain_3_reg ^ sbox_out_num_6_domain_4_reg ;



reg sbox_out_num_7_domain_1_reg,sbox_out_num_7_domain_2_reg,sbox_out_num_7_domain_3_reg,sbox_out_num_7_domain_4_reg ;
always@(posedge clk)
begin
	sbox_out_num_7_domain_1_reg <= inner_plus_cross_module_equation_num7_domain_1 ;
	sbox_out_num_7_domain_2_reg <= inner_plus_cross_module_equation_num7_domain_2 ^ rand_bit_second[8] ;
	sbox_out_num_7_domain_3_reg <= inner_plus_cross_module_equation_num7_domain_3 ^ rand_bit_second[8] ;
	sbox_out_num_7_domain_4_reg <= inner_plus_cross_module_equation_num7_domain_4 ;
end

wire sbox_out_num_7_share1, sbox_out_num_7_share2 ;
assign sbox_out_num_7_share1 = sbox_out_num_7_domain_1_reg ^ sbox_out_num_7_domain_2_reg ;
assign sbox_out_num_7_share2 = sbox_out_num_7_domain_3_reg ^ sbox_out_num_7_domain_4_reg ;



assign output_sbox_share1 = {sbox_out_num_7_share1,sbox_out_num_6_share1,sbox_out_num_5_share1,sbox_out_num_4_share1,sbox_out_num_3_share1,sbox_out_num_2_share1,sbox_out_num_1_share1,sbox_out_num_0_share1};
assign output_sbox_share2 = {sbox_out_num_7_share2,sbox_out_num_6_share2,sbox_out_num_5_share2,sbox_out_num_4_share2,sbox_out_num_3_share2,sbox_out_num_2_share2,sbox_out_num_1_share2,sbox_out_num_0_share2};

endmodule