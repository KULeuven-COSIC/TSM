`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: COSIC, KU Leuven, Belgium
// Engineer: Dilip Kumar S V
// Paper: Higher-Order Time Sharing Masking
// Authors: Dilip Kumar S. V., Siemen Dhooghe, Josep Balasch, Benedikt Gierlichs, Ingrid Verbauwhede
// Create Date: 22:00:00 02/22/2025
// Design Name: Combinatorial Logic for AES S-Box
// Module Name: combi_logic_cycle3_output_share2
// Project Name: AES Masked S-Box
// Target Device: FPGA
// Tool Versions: Vivado 2020.2
// Description: Contains combinatorial logic combining \( h_{\pi(I)} \) with \( g^2 \) functions 
//              to produce one share of the eight outputs of the AES S-box.
// Dependencies: None
//
// Revision:
// Revision 0.01 - Initial version
//
//////////////////////////////////////////////////////////////////////////////////

module combi_logic_cycle3_output_share2 (
    x0_subscript0_share2_reg , x2_subscript0_share2_reg , x3_subscript0_share2_reg , x4_subscript0_share2_reg , x6_subscript0_share2_reg , x7_subscript0_share2_reg , x1_subscript0_share2_reg , x5_subscript0_share2_reg , x0x1_subscript0_share2_reg , x0x4_subscript0_share2_reg , x0x5_subscript0_share2_reg , x0x6_subscript0_share2_reg , x1x2_subscript0_share2_reg , x1x3_subscript0_share2_reg , x1x4_subscript0_share2_reg , x1x6_subscript0_share2_reg , x2x3_subscript0_share2_reg , x2x4_subscript0_share2_reg , x2x6_subscript0_share2_reg , x2x7_subscript0_share2_reg , x4x6_subscript0_share2_reg , x5x6_subscript0_share2_reg , x5x7_subscript0_share2_reg , x6x7_subscript0_share2_reg , x0x2_subscript0_share2_reg , x0x3_subscript0_share2_reg , x0x7_subscript0_share2_reg , x1x7_subscript0_share2_reg , x3x7_subscript0_share2_reg , x4x5_subscript0_share2_reg , x3x4_subscript0_share2_reg , x4x7_subscript0_share2_reg , x3x6_subscript0_share2_reg , x1x5_subscript0_share2_reg , x2x5_subscript0_share2_reg , x3x5_subscript0_share2_reg , x0x1x4_subscript0_share2_reg , x0x1x6_subscript0_share2_reg , x0x1x7_subscript0_share2_reg , x0x2x4_subscript0_share2_reg , x0x2x5_subscript0_share2_reg , x0x2x6_subscript0_share2_reg , x0x2x7_subscript0_share2_reg , x0x3x4_subscript0_share2_reg , x0x3x5_subscript0_share2_reg , x0x3x6_subscript0_share2_reg , x0x4x6_subscript0_share2_reg , x0x4x7_subscript0_share2_reg , x1x2x3_subscript0_share2_reg , x1x2x4_subscript0_share2_reg , x1x2x6_subscript0_share2_reg , x1x3x4_subscript0_share2_reg , x1x3x7_subscript0_share2_reg , x1x4x6_subscript0_share2_reg , x1x5x6_subscript0_share2_reg , x2x3x5_subscript0_share2_reg , x2x3x7_subscript0_share2_reg , x2x4x7_subscript0_share2_reg , x2x5x6_subscript0_share2_reg , x2x5x7_subscript0_share2_reg , x2x6x7_subscript0_share2_reg , x3x4x7_subscript0_share2_reg , x3x5x7_subscript0_share2_reg , x3x6x7_subscript0_share2_reg , x4x5x6_subscript0_share2_reg , x5x6x7_subscript0_share2_reg , x0x1x3_subscript0_share2_reg , x0x2x3_subscript0_share2_reg , x0x4x5_subscript0_share2_reg , x0x5x7_subscript0_share2_reg , x0x6x7_subscript0_share2_reg , x1x3x5_subscript0_share2_reg , x1x3x6_subscript0_share2_reg , x1x4x7_subscript0_share2_reg , x2x3x4_subscript0_share2_reg , x2x3x6_subscript0_share2_reg , x3x4x6_subscript0_share2_reg , x3x5x6_subscript0_share2_reg , x0x1x5_subscript0_share2_reg , x0x3x7_subscript0_share2_reg , x1x2x5_subscript0_share2_reg , x1x2x7_subscript0_share2_reg , x1x4x5_subscript0_share2_reg , x1x5x7_subscript0_share2_reg , x2x4x5_subscript0_share2_reg , x3x4x5_subscript0_share2_reg , x4x6x7_subscript0_share2_reg , x1x6x7_subscript0_share2_reg , x4x5x7_subscript0_share2_reg , x0x1x2_subscript0_share2_reg , x0x5x6_subscript0_share2_reg , x2x4x6_subscript0_share2_reg , x0x1x2x3_subscript0_share2_reg , x0x1x2x5_subscript0_share2_reg , x0x1x2x6_subscript0_share2_reg , x0x1x2x7_subscript0_share2_reg , x0x1x4x5_subscript0_share2_reg , x0x1x4x7_subscript0_share2_reg , x0x2x3x5_subscript0_share2_reg , x0x2x3x7_subscript0_share2_reg , x0x2x4x5_subscript0_share2_reg , x0x2x4x7_subscript0_share2_reg , x0x2x5x6_subscript0_share2_reg , x0x2x5x7_subscript0_share2_reg , x0x3x4x6_subscript0_share2_reg , x0x3x5x6_subscript0_share2_reg , x0x4x5x6_subscript0_share2_reg , x0x4x5x7_subscript0_share2_reg , x0x4x6x7_subscript0_share2_reg , x1x2x3x5_subscript0_share2_reg , x1x2x3x6_subscript0_share2_reg , x1x2x3x7_subscript0_share2_reg , x1x2x4x6_subscript0_share2_reg , x1x2x4x7_subscript0_share2_reg , x1x2x6x7_subscript0_share2_reg , x1x3x4x6_subscript0_share2_reg , x1x3x6x7_subscript0_share2_reg , x1x4x5x6_subscript0_share2_reg , x1x4x5x7_subscript0_share2_reg , x1x5x6x7_subscript0_share2_reg , x2x3x5x7_subscript0_share2_reg , x2x3x6x7_subscript0_share2_reg , x2x4x5x6_subscript0_share2_reg , x2x4x5x7_subscript0_share2_reg , x3x5x6x7_subscript0_share2_reg , x0x1x3x4_subscript0_share2_reg , x0x1x3x6_subscript0_share2_reg , x0x1x5x6_subscript0_share2_reg , x0x2x3x6_subscript0_share2_reg , x0x3x4x5_subscript0_share2_reg , x1x2x5x6_subscript0_share2_reg , x1x2x5x7_subscript0_share2_reg , x1x3x4x5_subscript0_share2_reg , x1x3x4x7_subscript0_share2_reg , x1x3x5x6_subscript0_share2_reg , x1x3x5x7_subscript0_share2_reg , x1x4x6x7_subscript0_share2_reg , x2x3x4x5_subscript0_share2_reg , x2x3x4x7_subscript0_share2_reg , x2x4x6x7_subscript0_share2_reg , x3x4x5x6_subscript0_share2_reg , x3x4x5x7_subscript0_share2_reg , x3x4x6x7_subscript0_share2_reg , x0x1x3x5_subscript0_share2_reg , x0x1x4x6_subscript0_share2_reg , x0x2x3x4_subscript0_share2_reg , x0x2x4x6_subscript0_share2_reg , x0x3x4x7_subscript0_share2_reg , x0x3x5x7_subscript0_share2_reg , x1x2x3x4_subscript0_share2_reg , x2x3x4x6_subscript0_share2_reg , x2x3x5x6_subscript0_share2_reg , x2x5x6x7_subscript0_share2_reg , x4x5x6x7_subscript0_share2_reg , x0x1x2x4_subscript0_share2_reg , x0x1x6x7_subscript0_share2_reg , x0x2x6x7_subscript0_share2_reg , x0x3x6x7_subscript0_share2_reg , x0x5x6x7_subscript0_share2_reg , x1x2x4x5_subscript0_share2_reg , x0x1x3x7_subscript0_share2_reg , x0x1x5x7_subscript0_share2_reg , x0x1x2x3x4_subscript0_share2_reg , x0x1x2x3x6_subscript0_share2_reg , x0x1x2x3x7_subscript0_share2_reg , x0x1x2x4x5_subscript0_share2_reg , x0x1x2x4x7_subscript0_share2_reg , x0x1x2x5x7_subscript0_share2_reg , x0x1x2x6x7_subscript0_share2_reg , x0x1x3x4x6_subscript0_share2_reg , x0x1x3x5x6_subscript0_share2_reg , x0x1x3x5x7_subscript0_share2_reg , x0x1x3x6x7_subscript0_share2_reg , x0x1x4x5x6_subscript0_share2_reg , x0x1x5x6x7_subscript0_share2_reg , x0x2x3x4x5_subscript0_share2_reg , x0x2x3x4x6_subscript0_share2_reg , x0x2x4x5x7_subscript0_share2_reg , x0x2x4x6x7_subscript0_share2_reg , x0x3x4x5x6_subscript0_share2_reg , x0x3x4x5x7_subscript0_share2_reg , x0x3x4x6x7_subscript0_share2_reg , x0x3x5x6x7_subscript0_share2_reg , x1x2x3x5x6_subscript0_share2_reg , x1x2x3x5x7_subscript0_share2_reg , x1x2x4x5x6_subscript0_share2_reg , x1x2x4x6x7_subscript0_share2_reg , x1x2x5x6x7_subscript0_share2_reg , x1x3x4x5x7_subscript0_share2_reg , x2x3x4x5x6_subscript0_share2_reg , x2x3x4x5x7_subscript0_share2_reg , x2x4x5x6x7_subscript0_share2_reg , x0x1x2x4x6_subscript0_share2_reg , x0x1x3x4x7_subscript0_share2_reg , x0x2x3x4x7_subscript0_share2_reg , x0x2x3x5x7_subscript0_share2_reg , x0x2x3x6x7_subscript0_share2_reg , x0x2x4x5x6_subscript0_share2_reg , x0x2x5x6x7_subscript0_share2_reg , x0x4x5x6x7_subscript0_share2_reg , x1x2x3x4x6_subscript0_share2_reg , x1x3x4x5x6_subscript0_share2_reg , x2x3x4x6x7_subscript0_share2_reg , x0x1x2x3x5_subscript0_share2_reg , x0x1x4x6x7_subscript0_share2_reg , x1x2x3x4x5_subscript0_share2_reg , x1x2x3x6x7_subscript0_share2_reg , x1x2x4x5x7_subscript0_share2_reg , x1x3x4x6x7_subscript0_share2_reg , x1x3x5x6x7_subscript0_share2_reg , x1x4x5x6x7_subscript0_share2_reg , x2x3x5x6x7_subscript0_share2_reg , x3x4x5x6x7_subscript0_share2_reg , x0x1x2x5x6_subscript0_share2_reg , x0x1x3x4x5_subscript0_share2_reg , x0x1x4x5x7_subscript0_share2_reg , x0x2x3x5x6_subscript0_share2_reg , x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x4x6_subscript0_share2_reg , x0x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x5x7_subscript0_share2_reg , x0x1x2x3x6x7_subscript0_share2_reg , x0x1x2x4x5x7_subscript0_share2_reg , x0x1x2x5x6x7_subscript0_share2_reg , x0x1x3x4x6x7_subscript0_share2_reg , x0x1x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6_subscript0_share2_reg , x0x2x3x4x5x7_subscript0_share2_reg , x0x2x3x5x6x7_subscript0_share2_reg , x1x2x3x4x6x7_subscript0_share2_reg , x1x2x4x5x6x7_subscript0_share2_reg , x1x3x4x5x6x7_subscript0_share2_reg , x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6_subscript0_share2_reg , x0x1x2x4x6x7_subscript0_share2_reg , x0x1x3x4x5x6_subscript0_share2_reg , x0x2x3x4x6x7_subscript0_share2_reg , x1x2x3x4x5x6_subscript0_share2_reg , x1x2x3x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5_subscript0_share2_reg , x0x1x2x4x5x6_subscript0_share2_reg , x0x1x3x4x5x7_subscript0_share2_reg , x0x1x3x5x6x7_subscript0_share2_reg , x0x2x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x7_subscript0_share2_reg , x0x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x6x7_subscript0_share2_reg , x0x1x2x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6x7_subscript0_share2_reg , x0x1x3x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5x6_subscript0_share2_reg , x0x1x2x3x4x5x7_subscript0_share2_reg , 
    x0_share_in, x1_share_in, x2_share_in, x3_share_in, x4_share_in, x5_share_in, x6_share_in, x7_share_in ,
    sbox_out1_share2, sbox_out2_share2, sbox_out3_share2, sbox_out4_share2, sbox_out5_share2, sbox_out6_share2, sbox_out7_share2, sbox_out8_share2 
);

     
input  x0_subscript0_share2_reg , x2_subscript0_share2_reg , x3_subscript0_share2_reg , x4_subscript0_share2_reg , x6_subscript0_share2_reg , x7_subscript0_share2_reg , x1_subscript0_share2_reg , x5_subscript0_share2_reg , x0x1_subscript0_share2_reg , x0x4_subscript0_share2_reg , x0x5_subscript0_share2_reg , x0x6_subscript0_share2_reg , x1x2_subscript0_share2_reg , x1x3_subscript0_share2_reg , x1x4_subscript0_share2_reg , x1x6_subscript0_share2_reg , x2x3_subscript0_share2_reg , x2x4_subscript0_share2_reg , x2x6_subscript0_share2_reg , x2x7_subscript0_share2_reg , x4x6_subscript0_share2_reg , x5x6_subscript0_share2_reg , x5x7_subscript0_share2_reg , x6x7_subscript0_share2_reg , x0x2_subscript0_share2_reg , x0x3_subscript0_share2_reg , x0x7_subscript0_share2_reg , x1x7_subscript0_share2_reg , x3x7_subscript0_share2_reg , x4x5_subscript0_share2_reg , x3x4_subscript0_share2_reg , x4x7_subscript0_share2_reg , x3x6_subscript0_share2_reg , x1x5_subscript0_share2_reg , x2x5_subscript0_share2_reg , x3x5_subscript0_share2_reg , x0x1x4_subscript0_share2_reg , x0x1x6_subscript0_share2_reg , x0x1x7_subscript0_share2_reg , x0x2x4_subscript0_share2_reg , x0x2x5_subscript0_share2_reg , x0x2x6_subscript0_share2_reg , x0x2x7_subscript0_share2_reg , x0x3x4_subscript0_share2_reg , x0x3x5_subscript0_share2_reg , x0x3x6_subscript0_share2_reg , x0x4x6_subscript0_share2_reg , x0x4x7_subscript0_share2_reg , x1x2x3_subscript0_share2_reg , x1x2x4_subscript0_share2_reg , x1x2x6_subscript0_share2_reg , x1x3x4_subscript0_share2_reg , x1x3x7_subscript0_share2_reg , x1x4x6_subscript0_share2_reg , x1x5x6_subscript0_share2_reg , x2x3x5_subscript0_share2_reg , x2x3x7_subscript0_share2_reg , x2x4x7_subscript0_share2_reg , x2x5x6_subscript0_share2_reg , x2x5x7_subscript0_share2_reg , x2x6x7_subscript0_share2_reg , x3x4x7_subscript0_share2_reg , x3x5x7_subscript0_share2_reg , x3x6x7_subscript0_share2_reg , x4x5x6_subscript0_share2_reg , x5x6x7_subscript0_share2_reg , x0x1x3_subscript0_share2_reg , x0x2x3_subscript0_share2_reg , x0x4x5_subscript0_share2_reg , x0x5x7_subscript0_share2_reg , x0x6x7_subscript0_share2_reg , x1x3x5_subscript0_share2_reg , x1x3x6_subscript0_share2_reg , x1x4x7_subscript0_share2_reg , x2x3x4_subscript0_share2_reg , x2x3x6_subscript0_share2_reg , x3x4x6_subscript0_share2_reg , x3x5x6_subscript0_share2_reg , x0x1x5_subscript0_share2_reg , x0x3x7_subscript0_share2_reg , x1x2x5_subscript0_share2_reg , x1x2x7_subscript0_share2_reg , x1x4x5_subscript0_share2_reg , x1x5x7_subscript0_share2_reg , x2x4x5_subscript0_share2_reg , x3x4x5_subscript0_share2_reg , x4x6x7_subscript0_share2_reg , x1x6x7_subscript0_share2_reg , x4x5x7_subscript0_share2_reg , x0x1x2_subscript0_share2_reg , x0x5x6_subscript0_share2_reg , x2x4x6_subscript0_share2_reg , x0x1x2x3_subscript0_share2_reg , x0x1x2x5_subscript0_share2_reg , x0x1x2x6_subscript0_share2_reg , x0x1x2x7_subscript0_share2_reg , x0x1x4x5_subscript0_share2_reg , x0x1x4x7_subscript0_share2_reg , x0x2x3x5_subscript0_share2_reg , x0x2x3x7_subscript0_share2_reg , x0x2x4x5_subscript0_share2_reg , x0x2x4x7_subscript0_share2_reg , x0x2x5x6_subscript0_share2_reg , x0x2x5x7_subscript0_share2_reg , x0x3x4x6_subscript0_share2_reg , x0x3x5x6_subscript0_share2_reg , x0x4x5x6_subscript0_share2_reg , x0x4x5x7_subscript0_share2_reg , x0x4x6x7_subscript0_share2_reg , x1x2x3x5_subscript0_share2_reg , x1x2x3x6_subscript0_share2_reg , x1x2x3x7_subscript0_share2_reg , x1x2x4x6_subscript0_share2_reg , x1x2x4x7_subscript0_share2_reg , x1x2x6x7_subscript0_share2_reg , x1x3x4x6_subscript0_share2_reg , x1x3x6x7_subscript0_share2_reg , x1x4x5x6_subscript0_share2_reg , x1x4x5x7_subscript0_share2_reg , x1x5x6x7_subscript0_share2_reg , x2x3x5x7_subscript0_share2_reg , x2x3x6x7_subscript0_share2_reg , x2x4x5x6_subscript0_share2_reg , x2x4x5x7_subscript0_share2_reg , x3x5x6x7_subscript0_share2_reg , x0x1x3x4_subscript0_share2_reg , x0x1x3x6_subscript0_share2_reg , x0x1x5x6_subscript0_share2_reg , x0x2x3x6_subscript0_share2_reg , x0x3x4x5_subscript0_share2_reg , x1x2x5x6_subscript0_share2_reg , x1x2x5x7_subscript0_share2_reg , x1x3x4x5_subscript0_share2_reg , x1x3x4x7_subscript0_share2_reg , x1x3x5x6_subscript0_share2_reg , x1x3x5x7_subscript0_share2_reg , x1x4x6x7_subscript0_share2_reg , x2x3x4x5_subscript0_share2_reg , x2x3x4x7_subscript0_share2_reg , x2x4x6x7_subscript0_share2_reg , x3x4x5x6_subscript0_share2_reg , x3x4x5x7_subscript0_share2_reg , x3x4x6x7_subscript0_share2_reg , x0x1x3x5_subscript0_share2_reg , x0x1x4x6_subscript0_share2_reg , x0x2x3x4_subscript0_share2_reg , x0x2x4x6_subscript0_share2_reg , x0x3x4x7_subscript0_share2_reg , x0x3x5x7_subscript0_share2_reg , x1x2x3x4_subscript0_share2_reg , x2x3x4x6_subscript0_share2_reg , x2x3x5x6_subscript0_share2_reg , x2x5x6x7_subscript0_share2_reg , x4x5x6x7_subscript0_share2_reg , x0x1x2x4_subscript0_share2_reg , x0x1x6x7_subscript0_share2_reg , x0x2x6x7_subscript0_share2_reg , x0x3x6x7_subscript0_share2_reg , x0x5x6x7_subscript0_share2_reg , x1x2x4x5_subscript0_share2_reg , x0x1x3x7_subscript0_share2_reg , x0x1x5x7_subscript0_share2_reg , x0x1x2x3x4_subscript0_share2_reg , x0x1x2x3x6_subscript0_share2_reg , x0x1x2x3x7_subscript0_share2_reg , x0x1x2x4x5_subscript0_share2_reg , x0x1x2x4x7_subscript0_share2_reg , x0x1x2x5x7_subscript0_share2_reg , x0x1x2x6x7_subscript0_share2_reg , x0x1x3x4x6_subscript0_share2_reg , x0x1x3x5x6_subscript0_share2_reg , x0x1x3x5x7_subscript0_share2_reg , x0x1x3x6x7_subscript0_share2_reg , x0x1x4x5x6_subscript0_share2_reg , x0x1x5x6x7_subscript0_share2_reg , x0x2x3x4x5_subscript0_share2_reg , x0x2x3x4x6_subscript0_share2_reg , x0x2x4x5x7_subscript0_share2_reg , x0x2x4x6x7_subscript0_share2_reg , x0x3x4x5x6_subscript0_share2_reg , x0x3x4x5x7_subscript0_share2_reg , x0x3x4x6x7_subscript0_share2_reg , x0x3x5x6x7_subscript0_share2_reg , x1x2x3x5x6_subscript0_share2_reg , x1x2x3x5x7_subscript0_share2_reg , x1x2x4x5x6_subscript0_share2_reg , x1x2x4x6x7_subscript0_share2_reg , x1x2x5x6x7_subscript0_share2_reg , x1x3x4x5x7_subscript0_share2_reg , x2x3x4x5x6_subscript0_share2_reg , x2x3x4x5x7_subscript0_share2_reg , x2x4x5x6x7_subscript0_share2_reg , x0x1x2x4x6_subscript0_share2_reg , x0x1x3x4x7_subscript0_share2_reg , x0x2x3x4x7_subscript0_share2_reg , x0x2x3x5x7_subscript0_share2_reg , x0x2x3x6x7_subscript0_share2_reg , x0x2x4x5x6_subscript0_share2_reg , x0x2x5x6x7_subscript0_share2_reg , x0x4x5x6x7_subscript0_share2_reg , x1x2x3x4x6_subscript0_share2_reg , x1x3x4x5x6_subscript0_share2_reg , x2x3x4x6x7_subscript0_share2_reg , x0x1x2x3x5_subscript0_share2_reg , x0x1x4x6x7_subscript0_share2_reg , x1x2x3x4x5_subscript0_share2_reg , x1x2x3x6x7_subscript0_share2_reg , x1x2x4x5x7_subscript0_share2_reg , x1x3x4x6x7_subscript0_share2_reg , x1x3x5x6x7_subscript0_share2_reg , x1x4x5x6x7_subscript0_share2_reg , x2x3x5x6x7_subscript0_share2_reg , x3x4x5x6x7_subscript0_share2_reg , x0x1x2x5x6_subscript0_share2_reg , x0x1x3x4x5_subscript0_share2_reg , x0x1x4x5x7_subscript0_share2_reg , x0x2x3x5x6_subscript0_share2_reg , x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x4x6_subscript0_share2_reg , x0x1x2x3x4x7_subscript0_share2_reg , x0x1x2x3x5x7_subscript0_share2_reg , x0x1x2x3x6x7_subscript0_share2_reg , x0x1x2x4x5x7_subscript0_share2_reg , x0x1x2x5x6x7_subscript0_share2_reg , x0x1x3x4x6x7_subscript0_share2_reg , x0x1x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6_subscript0_share2_reg , x0x2x3x4x5x7_subscript0_share2_reg , x0x2x3x5x6x7_subscript0_share2_reg , x1x2x3x4x6x7_subscript0_share2_reg , x1x2x4x5x6x7_subscript0_share2_reg , x1x3x4x5x6x7_subscript0_share2_reg , x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6_subscript0_share2_reg , x0x1x2x4x6x7_subscript0_share2_reg , x0x1x3x4x5x6_subscript0_share2_reg , x0x2x3x4x6x7_subscript0_share2_reg , x1x2x3x4x5x6_subscript0_share2_reg , x1x2x3x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5_subscript0_share2_reg , x0x1x2x4x5x6_subscript0_share2_reg , x0x1x3x4x5x7_subscript0_share2_reg , x0x1x3x5x6x7_subscript0_share2_reg , x0x2x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x7_subscript0_share2_reg , x0x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x6x7_subscript0_share2_reg , x0x1x2x4x5x6x7_subscript0_share2_reg , x0x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x5x6x7_subscript0_share2_reg , x0x1x3x4x5x6x7_subscript0_share2_reg , x1x2x3x4x5x6x7_subscript0_share2_reg , x0x1x2x3x4x5x6_subscript0_share2_reg , x0x1x2x3x4x5x7_subscript0_share2_reg ;
input  x0_share_in, x1_share_in, x2_share_in, x3_share_in, x4_share_in, x5_share_in, x6_share_in, x7_share_in ;


output sbox_out1_share2, sbox_out2_share2, sbox_out3_share2, sbox_out4_share2, sbox_out5_share2, sbox_out6_share2, sbox_out7_share2, sbox_out8_share2 ;

wire x0_second_share, x1_second_share, x2_second_share, x3_second_share, x4_second_share, x5_second_share, x6_second_share, x7_second_share ;
wire x0x1_second_share , x0x2_second_share , x0x3_second_share , x0x4_second_share , x0x5_second_share , x0x6_second_share , x0x7_second_share , x1x2_second_share , x1x3_second_share , x1x4_second_share , x1x5_second_share , x1x6_second_share , x1x7_second_share , x2x3_second_share , x2x4_second_share , x2x5_second_share , x2x6_second_share , x2x7_second_share , x3x4_second_share , x3x5_second_share , x3x6_second_share , x3x7_second_share , x4x5_second_share , x4x6_second_share , x4x7_second_share , x5x6_second_share , x5x7_second_share , x6x7_second_share , x0x1x2_second_share , x0x1x3_second_share , x0x1x4_second_share , x0x1x5_second_share , x0x1x6_second_share , x0x1x7_second_share , x0x2x3_second_share , x0x2x4_second_share , x0x2x5_second_share , x0x2x6_second_share , x0x2x7_second_share , x0x3x4_second_share , x0x3x5_second_share , x0x3x6_second_share , x0x3x7_second_share , x0x4x5_second_share , x0x4x6_second_share , x0x4x7_second_share , x0x5x6_second_share , x0x5x7_second_share , x0x6x7_second_share , x1x2x3_second_share , x1x2x4_second_share , x1x2x5_second_share , x1x2x6_second_share , x1x2x7_second_share , x1x3x4_second_share , x1x3x5_second_share , x1x3x6_second_share , x1x3x7_second_share , x1x4x5_second_share , x1x4x6_second_share , x1x4x7_second_share , x1x5x6_second_share , x1x5x7_second_share , x1x6x7_second_share , x2x3x4_second_share , x2x3x5_second_share , x2x3x6_second_share , x2x3x7_second_share , x2x4x5_second_share , x2x4x6_second_share , x2x4x7_second_share , x2x5x6_second_share , x2x5x7_second_share , x2x6x7_second_share , x3x4x5_second_share , x3x4x6_second_share , x3x4x7_second_share , x3x5x6_second_share , x3x5x7_second_share , x3x6x7_second_share , x4x5x6_second_share , x4x5x7_second_share , x4x6x7_second_share , x5x6x7_second_share , x0x1x2x3_second_share , x0x1x2x4_second_share , x0x1x2x5_second_share , x0x1x2x6_second_share , x0x1x2x7_second_share , x0x1x3x4_second_share , x0x1x3x5_second_share , x0x1x3x6_second_share , x0x1x3x7_second_share , x0x1x4x5_second_share , x0x1x4x6_second_share , x0x1x4x7_second_share , x0x1x5x6_second_share , x0x1x5x7_second_share , x0x1x6x7_second_share , x0x2x3x4_second_share , x0x2x3x5_second_share , x0x2x3x6_second_share , x0x2x3x7_second_share , x0x2x4x5_second_share , x0x2x4x6_second_share , x0x2x4x7_second_share , x0x2x5x6_second_share , x0x2x5x7_second_share , x0x2x6x7_second_share , x0x3x4x5_second_share , x0x3x4x6_second_share , x0x3x4x7_second_share , x0x3x5x6_second_share , x0x3x5x7_second_share , x0x3x6x7_second_share , x0x4x5x6_second_share , x0x4x5x7_second_share , x0x4x6x7_second_share , x0x5x6x7_second_share , x1x2x3x4_second_share , x1x2x3x5_second_share , x1x2x3x6_second_share , x1x2x3x7_second_share , x1x2x4x5_second_share , x1x2x4x6_second_share , x1x2x4x7_second_share , x1x2x5x6_second_share , x1x2x5x7_second_share , x1x2x6x7_second_share , x1x3x4x5_second_share , x1x3x4x6_second_share , x1x3x4x7_second_share , x1x3x5x6_second_share , x1x3x5x7_second_share , x1x3x6x7_second_share , x1x4x5x6_second_share , x1x4x5x7_second_share , x1x4x6x7_second_share , x1x5x6x7_second_share , x2x3x4x5_second_share , x2x3x4x6_second_share , x2x3x4x7_second_share , x2x3x5x6_second_share , x2x3x5x7_second_share , x2x3x6x7_second_share , x2x4x5x6_second_share , x2x4x5x7_second_share , x2x4x6x7_second_share , x2x5x6x7_second_share , x3x4x5x6_second_share , x3x4x5x7_second_share , x3x4x6x7_second_share , x3x5x6x7_second_share , x4x5x6x7_second_share , x0x1x2x3x4_second_share , x0x1x2x3x5_second_share , x0x1x2x3x6_second_share , x0x1x2x3x7_second_share , x0x1x2x4x5_second_share , x0x1x2x4x6_second_share , x0x1x2x4x7_second_share , x0x1x2x5x6_second_share , x0x1x2x5x7_second_share , x0x1x2x6x7_second_share , x0x1x3x4x5_second_share , x0x1x3x4x6_second_share , x0x1x3x4x7_second_share , x0x1x3x5x6_second_share , x0x1x3x5x7_second_share , x0x1x3x6x7_second_share , x0x1x4x5x6_second_share , x0x1x4x5x7_second_share , x0x1x4x6x7_second_share , x0x1x5x6x7_second_share , x0x2x3x4x5_second_share , x0x2x3x4x6_second_share , x0x2x3x4x7_second_share , x0x2x3x5x6_second_share , x0x2x3x5x7_second_share , x0x2x3x6x7_second_share , x0x2x4x5x6_second_share , x0x2x4x5x7_second_share , x0x2x4x6x7_second_share , x0x2x5x6x7_second_share , x0x3x4x5x6_second_share , x0x3x4x5x7_second_share , x0x3x4x6x7_second_share , x0x3x5x6x7_second_share , x0x4x5x6x7_second_share , x1x2x3x4x5_second_share , x1x2x3x4x6_second_share , x1x2x3x4x7_second_share , x1x2x3x5x6_second_share , x1x2x3x5x7_second_share , x1x2x3x6x7_second_share , x1x2x4x5x6_second_share , x1x2x4x5x7_second_share , x1x2x4x6x7_second_share , x1x2x5x6x7_second_share , x1x3x4x5x6_second_share , x1x3x4x5x7_second_share , x1x3x4x6x7_second_share , x1x3x5x6x7_second_share , x1x4x5x6x7_second_share , x2x3x4x5x6_second_share , x2x3x4x5x7_second_share , x2x3x4x6x7_second_share , x2x3x5x6x7_second_share , x2x4x5x6x7_second_share , x3x4x5x6x7_second_share , x0x1x2x3x4x5_second_share , x0x1x2x3x4x6_second_share , x0x1x2x3x4x7_second_share , x0x1x2x3x5x6_second_share , x0x1x2x3x5x7_second_share , x0x1x2x3x6x7_second_share , x0x1x2x4x5x6_second_share , x0x1x2x4x5x7_second_share , x0x1x2x4x6x7_second_share , x0x1x2x5x6x7_second_share , x0x1x3x4x5x6_second_share , x0x1x3x4x5x7_second_share , x0x1x3x4x6x7_second_share , x0x1x3x5x6x7_second_share , x0x1x4x5x6x7_second_share , x0x2x3x4x5x6_second_share , x0x2x3x4x5x7_second_share , x0x2x3x4x6x7_second_share , x0x2x3x5x6x7_second_share , x0x2x4x5x6x7_second_share , x0x3x4x5x6x7_second_share , x1x2x3x4x5x6_second_share , x1x2x3x4x5x7_second_share , x1x2x3x4x6x7_second_share , x1x2x3x5x6x7_second_share , x1x2x4x5x6x7_second_share , x1x3x4x5x6x7_second_share , x2x3x4x5x6x7_second_share , x0x1x2x3x4x5x6_second_share , x0x1x2x3x4x5x7_second_share , x0x1x2x3x4x6x7_second_share , x0x1x2x3x5x6x7_second_share , x0x1x2x4x5x6x7_second_share , x0x1x3x4x5x6x7_second_share , x0x2x3x4x5x6x7_second_share , x1x2x3x4x5x6x7_second_share ;

// All crossproducts

assign x0_share2_reg             =  x0_share_in ;
assign x1_share2_reg             =  x1_share_in ;
assign x2_share2_reg             =  x2_share_in ;
assign x3_share2_reg             =  x3_share_in ;
assign x4_share2_reg             =  x4_share_in ;
assign x5_share2_reg             =  x5_share_in ;
assign x6_share2_reg             =  x6_share_in ;
assign x7_share2_reg             =  x7_share_in ;
assign x0x1_share2_reg           =  x0_share_in & x1_share_in   ;
assign x0x4_share2_reg           =  x0_share_in & x4_share_in   ;
assign x0x5_share2_reg           =  x0_share_in & x5_share_in   ;
assign x0x6_share2_reg           =  x0_share_in & x6_share_in   ;
assign x1x2_share2_reg           =  x1_share_in & x2_share_in   ;
assign x1x3_share2_reg           =  x1_share_in & x3_share_in   ;
assign x1x4_share2_reg           =  x1_share_in & x4_share_in   ;
assign x1x6_share2_reg           =  x1_share_in & x6_share_in   ;
assign x2x3_share2_reg           =  x2_share_in & x3_share_in   ;
assign x2x4_share2_reg           =  x2_share_in & x4_share_in   ;
assign x2x6_share2_reg           =  x2_share_in & x6_share_in   ;
assign x2x7_share2_reg           =  x2_share_in & x7_share_in   ;
assign x4x6_share2_reg           =  x4_share_in & x6_share_in   ;
assign x5x6_share2_reg           =  x5_share_in & x6_share_in   ;
assign x5x7_share2_reg           =  x5_share_in & x7_share_in   ;
assign x6x7_share2_reg           =  x6_share_in & x7_share_in   ;
assign x0x2_share2_reg           =  x0_share_in & x2_share_in   ;
assign x0x3_share2_reg           =  x0_share_in & x3_share_in   ;
assign x0x7_share2_reg           =  x0_share_in & x7_share_in   ;
assign x1x7_share2_reg           =  x1_share_in & x7_share_in   ;
assign x3x7_share2_reg           =  x3_share_in & x7_share_in   ;
assign x4x5_share2_reg           =  x4_share_in & x5_share_in   ;
assign x3x4_share2_reg           =  x3_share_in & x4_share_in   ;
assign x4x7_share2_reg           =  x4_share_in & x7_share_in   ;
assign x3x6_share2_reg           =  x3_share_in & x6_share_in   ;
assign x1x5_share2_reg           =  x1_share_in & x5_share_in   ;
assign x2x5_share2_reg           =  x2_share_in & x5_share_in   ;
assign x3x5_share2_reg           =  x3_share_in & x5_share_in   ;
assign x0x1x4_share2_reg         =  x0_share_in & x1_share_in & x4_share_in   ;
assign x0x1x6_share2_reg         =  x0_share_in & x1_share_in & x6_share_in   ;
assign x0x1x7_share2_reg         =  x0_share_in & x1_share_in & x7_share_in   ;
assign x0x2x4_share2_reg         =  x0_share_in & x2_share_in & x4_share_in   ;
assign x0x2x5_share2_reg         =  x0_share_in & x2_share_in & x5_share_in   ;
assign x0x2x6_share2_reg         =  x0_share_in & x2_share_in & x6_share_in   ;
assign x0x2x7_share2_reg         =  x0_share_in & x2_share_in & x7_share_in   ;
assign x0x3x4_share2_reg         =  x0_share_in & x3_share_in & x4_share_in   ;
assign x0x3x5_share2_reg         =  x0_share_in & x3_share_in & x5_share_in   ;
assign x0x3x6_share2_reg         =  x0_share_in & x3_share_in & x6_share_in   ;
assign x0x4x6_share2_reg         =  x0_share_in & x4_share_in & x6_share_in   ;
assign x0x4x7_share2_reg         =  x0_share_in & x4_share_in & x7_share_in   ;
assign x1x2x3_share2_reg         =  x1_share_in & x2_share_in & x3_share_in   ;
assign x1x2x4_share2_reg         =  x1_share_in & x2_share_in & x4_share_in   ;
assign x1x2x6_share2_reg         =  x1_share_in & x2_share_in & x6_share_in   ;
assign x1x3x4_share2_reg         =  x1_share_in & x3_share_in & x4_share_in   ;
assign x1x3x7_share2_reg         =  x1_share_in & x3_share_in & x7_share_in   ;
assign x1x4x6_share2_reg         =  x1_share_in & x4_share_in & x6_share_in   ;
assign x1x5x6_share2_reg         =  x1_share_in & x5_share_in & x6_share_in   ;
assign x2x3x5_share2_reg         =  x2_share_in & x3_share_in & x5_share_in   ;
assign x2x3x7_share2_reg         =  x2_share_in & x3_share_in & x7_share_in   ;
assign x2x4x7_share2_reg         =  x2_share_in & x4_share_in & x7_share_in   ;
assign x2x5x6_share2_reg         =  x2_share_in & x5_share_in & x6_share_in   ;
assign x2x5x7_share2_reg         =  x2_share_in & x5_share_in & x7_share_in   ;
assign x2x6x7_share2_reg         =  x2_share_in & x6_share_in & x7_share_in   ;
assign x3x4x7_share2_reg         =  x3_share_in & x4_share_in & x7_share_in   ;
assign x3x5x7_share2_reg         =  x3_share_in & x5_share_in & x7_share_in   ;
assign x3x6x7_share2_reg         =  x3_share_in & x6_share_in & x7_share_in   ;
assign x4x5x6_share2_reg         =  x4_share_in & x5_share_in & x6_share_in   ;
assign x5x6x7_share2_reg         =  x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3_share2_reg         =  x0_share_in & x1_share_in & x3_share_in   ;
assign x0x2x3_share2_reg         =  x0_share_in & x2_share_in & x3_share_in   ;
assign x0x4x5_share2_reg         =  x0_share_in & x4_share_in & x5_share_in   ;
assign x0x5x7_share2_reg         =  x0_share_in & x5_share_in & x7_share_in   ;
assign x0x6x7_share2_reg         =  x0_share_in & x6_share_in & x7_share_in   ;
assign x1x3x5_share2_reg         =  x1_share_in & x3_share_in & x5_share_in   ;
assign x1x3x6_share2_reg         =  x1_share_in & x3_share_in & x6_share_in   ;
assign x1x4x7_share2_reg         =  x1_share_in & x4_share_in & x7_share_in   ;
assign x2x3x4_share2_reg         =  x2_share_in & x3_share_in & x4_share_in   ;
assign x2x3x6_share2_reg         =  x2_share_in & x3_share_in & x6_share_in   ;
assign x3x4x6_share2_reg         =  x3_share_in & x4_share_in & x6_share_in   ;
assign x3x5x6_share2_reg         =  x3_share_in & x5_share_in & x6_share_in   ;
assign x0x1x5_share2_reg         =  x0_share_in & x1_share_in & x5_share_in   ;
assign x0x3x7_share2_reg         =  x0_share_in & x3_share_in & x7_share_in   ;
assign x1x2x5_share2_reg         =  x1_share_in & x2_share_in & x5_share_in   ;
assign x1x2x7_share2_reg         =  x1_share_in & x2_share_in & x7_share_in   ;
assign x1x4x5_share2_reg         =  x1_share_in & x4_share_in & x5_share_in   ;
assign x1x5x7_share2_reg         =  x1_share_in & x5_share_in & x7_share_in   ;
assign x2x4x5_share2_reg         =  x2_share_in & x4_share_in & x5_share_in   ;
assign x3x4x5_share2_reg         =  x3_share_in & x4_share_in & x5_share_in   ;
assign x4x6x7_share2_reg         =  x4_share_in & x6_share_in & x7_share_in   ;
assign x1x6x7_share2_reg         =  x1_share_in & x6_share_in & x7_share_in   ;
assign x4x5x7_share2_reg         =  x4_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2_share2_reg         =  x0_share_in & x1_share_in & x2_share_in   ;
assign x0x5x6_share2_reg         =  x0_share_in & x5_share_in & x6_share_in   ;
assign x2x4x6_share2_reg         =  x2_share_in & x4_share_in & x6_share_in   ;
assign x0x1x2x3_share2_reg       =  x0_share_in & x1_share_in & x2_share_in & x3_share_in   ;
assign x0x1x2x5_share2_reg       =  x0_share_in & x1_share_in & x2_share_in & x5_share_in   ;
assign x0x1x2x6_share2_reg       =  x0_share_in & x1_share_in & x2_share_in & x6_share_in   ;
assign x0x1x2x7_share2_reg       =  x0_share_in & x1_share_in & x2_share_in & x7_share_in   ;
assign x0x1x4x5_share2_reg       =  x0_share_in & x1_share_in & x4_share_in & x5_share_in   ;
assign x0x1x4x7_share2_reg       =  x0_share_in & x1_share_in & x4_share_in & x7_share_in   ;
assign x0x2x3x5_share2_reg       =  x0_share_in & x2_share_in & x3_share_in & x5_share_in   ;
assign x0x2x3x7_share2_reg       =  x0_share_in & x2_share_in & x3_share_in & x7_share_in   ;
assign x0x2x4x5_share2_reg       =  x0_share_in & x2_share_in & x4_share_in & x5_share_in   ;
assign x0x2x4x7_share2_reg       =  x0_share_in & x2_share_in & x4_share_in & x7_share_in   ;
assign x0x2x5x6_share2_reg       =  x0_share_in & x2_share_in & x5_share_in & x6_share_in   ;
assign x0x2x5x7_share2_reg       =  x0_share_in & x2_share_in & x5_share_in & x7_share_in   ;
assign x0x3x4x6_share2_reg       =  x0_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x0x3x5x6_share2_reg       =  x0_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x0x4x5x6_share2_reg       =  x0_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x4x5x7_share2_reg       =  x0_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x4x6x7_share2_reg       =  x0_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x5_share2_reg       =  x1_share_in & x2_share_in & x3_share_in & x5_share_in   ;
assign x1x2x3x6_share2_reg       =  x1_share_in & x2_share_in & x3_share_in & x6_share_in   ;
assign x1x2x3x7_share2_reg       =  x1_share_in & x2_share_in & x3_share_in & x7_share_in   ;
assign x1x2x4x6_share2_reg       =  x1_share_in & x2_share_in & x4_share_in & x6_share_in   ;
assign x1x2x4x7_share2_reg       =  x1_share_in & x2_share_in & x4_share_in & x7_share_in   ;
assign x1x2x6x7_share2_reg       =  x1_share_in & x2_share_in & x6_share_in & x7_share_in   ;
assign x1x3x4x6_share2_reg       =  x1_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x1x3x6x7_share2_reg       =  x1_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x1x4x5x6_share2_reg       =  x1_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x1x4x5x7_share2_reg       =  x1_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x1x5x6x7_share2_reg       =  x1_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x2x3x5x7_share2_reg       =  x2_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x2x3x6x7_share2_reg       =  x2_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x2x4x5x6_share2_reg       =  x2_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x2x4x5x7_share2_reg       =  x2_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x3x5x6x7_share2_reg       =  x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4_share2_reg       =  x0_share_in & x1_share_in & x3_share_in & x4_share_in   ;
assign x0x1x3x6_share2_reg       =  x0_share_in & x1_share_in & x3_share_in & x6_share_in   ;
assign x0x1x5x6_share2_reg       =  x0_share_in & x1_share_in & x5_share_in & x6_share_in   ;
assign x0x2x3x6_share2_reg       =  x0_share_in & x2_share_in & x3_share_in & x6_share_in   ;
assign x0x3x4x5_share2_reg       =  x0_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x1x2x5x6_share2_reg       =  x1_share_in & x2_share_in & x5_share_in & x6_share_in   ;
assign x1x2x5x7_share2_reg       =  x1_share_in & x2_share_in & x5_share_in & x7_share_in   ;
assign x1x3x4x5_share2_reg       =  x1_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x1x3x4x7_share2_reg       =  x1_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x1x3x5x6_share2_reg       =  x1_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x1x3x5x7_share2_reg       =  x1_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x1x4x6x7_share2_reg       =  x1_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x2x3x4x5_share2_reg       =  x2_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x2x3x4x7_share2_reg       =  x2_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x2x4x6x7_share2_reg       =  x2_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x3x4x5x6_share2_reg       =  x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x3x4x5x7_share2_reg       =  x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x3x4x6x7_share2_reg       =  x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x5_share2_reg       =  x0_share_in & x1_share_in & x3_share_in & x5_share_in   ;
assign x0x1x4x6_share2_reg       =  x0_share_in & x1_share_in & x4_share_in & x6_share_in   ;
assign x0x2x3x4_share2_reg       =  x0_share_in & x2_share_in & x3_share_in & x4_share_in   ;
assign x0x2x4x6_share2_reg       =  x0_share_in & x2_share_in & x4_share_in & x6_share_in   ;
assign x0x3x4x7_share2_reg       =  x0_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x3x5x7_share2_reg       =  x0_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x1x2x3x4_share2_reg       =  x1_share_in & x2_share_in & x3_share_in & x4_share_in   ;
assign x2x3x4x6_share2_reg       =  x2_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x2x3x5x6_share2_reg       =  x2_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x2x5x6x7_share2_reg       =  x2_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x4x5x6x7_share2_reg       =  x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x4_share2_reg       =  x0_share_in & x1_share_in & x2_share_in & x4_share_in   ;
assign x0x1x6x7_share2_reg       =  x0_share_in & x1_share_in & x6_share_in & x7_share_in   ;
assign x0x2x6x7_share2_reg       =  x0_share_in & x2_share_in & x6_share_in & x7_share_in   ;
assign x0x3x6x7_share2_reg       =  x0_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x0x5x6x7_share2_reg       =  x0_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x4x5_share2_reg       =  x1_share_in & x2_share_in & x4_share_in & x5_share_in   ;
assign x0x1x3x7_share2_reg       =  x0_share_in & x1_share_in & x3_share_in & x7_share_in   ;
assign x0x1x5x7_share2_reg       =  x0_share_in & x1_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2x3x4_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in   ;
assign x0x1x2x3x6_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x6_share_in   ;
assign x0x1x2x3x7_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x7_share_in   ;
assign x0x1x2x4x5_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x5_share_in   ;
assign x0x1x2x4x7_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x7_share_in   ;
assign x0x1x2x5x7_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2x6x7_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4x6_share2_reg     =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x0x1x3x5x6_share2_reg     =  x0_share_in & x1_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x0x1x3x5x7_share2_reg     =  x0_share_in & x1_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x0x1x3x6x7_share2_reg     =  x0_share_in & x1_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x0x1x4x5x6_share2_reg     =  x0_share_in & x1_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x1x5x6x7_share2_reg     =  x0_share_in & x1_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x2x3x4x5_share2_reg     =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x0x2x3x4x6_share2_reg     =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x0x2x4x5x7_share2_reg     =  x0_share_in & x2_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x2x4x6x7_share2_reg     =  x0_share_in & x2_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x3x4x5x6_share2_reg     =  x0_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x3x4x5x7_share2_reg     =  x0_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x3x4x6x7_share2_reg     =  x0_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x3x5x6x7_share2_reg     =  x0_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x5x6_share2_reg     =  x1_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x1x2x3x5x7_share2_reg     =  x1_share_in & x2_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x1x2x4x5x6_share2_reg     =  x1_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x1x2x4x6x7_share2_reg     =  x1_share_in & x2_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x5x6x7_share2_reg     =  x1_share_in & x2_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x3x4x5x7_share2_reg     =  x1_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x2x3x4x5x6_share2_reg     =  x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x2x3x4x5x7_share2_reg     =  x2_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x2x4x5x6x7_share2_reg     =  x2_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x4x6_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x6_share_in   ;
assign x0x1x3x4x7_share2_reg     =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x2x3x4x7_share2_reg     =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x2x3x5x7_share2_reg     =  x0_share_in & x2_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x0x2x3x6x7_share2_reg     =  x0_share_in & x2_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x0x2x4x5x6_share2_reg     =  x0_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x2x5x6x7_share2_reg     =  x0_share_in & x2_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x4x5x6x7_share2_reg     =  x0_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x6_share2_reg     =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x1x3x4x5x6_share2_reg     =  x1_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x2x3x4x6x7_share2_reg     =  x2_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x5_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x5_share_in   ;
assign x0x1x4x6x7_share2_reg     =  x0_share_in & x1_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x5_share2_reg     =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x1x2x3x6x7_share2_reg     =  x1_share_in & x2_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x1x2x4x5x7_share2_reg     =  x1_share_in & x2_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x1x3x4x6x7_share2_reg     =  x1_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x3x5x6x7_share2_reg     =  x1_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x4x5x6x7_share2_reg     =  x1_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x2x3x5x6x7_share2_reg     =  x2_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x3x4x5x6x7_share2_reg     =  x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x5x6_share2_reg     =  x0_share_in & x1_share_in & x2_share_in & x5_share_in & x6_share_in   ;
assign x0x1x3x4x5_share2_reg     =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x0x1x4x5x7_share2_reg     =  x0_share_in & x1_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x2x3x5x6_share2_reg     =  x0_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x1x2x3x4x7_share2_reg     =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x1x2x3x4x6_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in   ;
assign x0x1x2x3x4x7_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x7_share_in   ;
assign x0x1x2x3x5x7_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2x3x6x7_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x4x5x7_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x1x2x5x6x7_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4x6x7_share2_reg   =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x4x5x6x7_share2_reg   =  x0_share_in & x1_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x2x3x4x5x6_share2_reg   =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x2x3x4x5x7_share2_reg   =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x2x3x5x6x7_share2_reg   =  x0_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x6x7_share2_reg   =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x4x5x6x7_share2_reg   =  x1_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x3x4x5x6x7_share2_reg   =  x1_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x2x3x4x5x6x7_share2_reg   =  x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x5x6_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in   ;
assign x0x1x2x4x6x7_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4x5x6_share2_reg   =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x2x3x4x6x7_share2_reg   =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x5x6_share2_reg   =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x1x2x3x5x6x7_share2_reg   =  x1_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x4x5_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in   ;
assign x0x1x2x4x5x6_share2_reg   =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x1x3x4x5x7_share2_reg   =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x1x3x5x6x7_share2_reg   =  x0_share_in & x1_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x2x4x5x6x7_share2_reg   =  x0_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x5x7_share2_reg   =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;
assign x0x3x4x5x6x7_share2_reg   =  x0_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x4x6x7_share2_reg =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x4x5x6x7_share2_reg =  x0_share_in & x1_share_in & x2_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x2x3x4x5x6x7_share2_reg =  x0_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x5x6x7_share2_reg =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x3x4x5x6x7_share2_reg =  x0_share_in & x1_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x1x2x3x4x5x6x7_share2_reg =  x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in & x7_share_in   ;
assign x0x1x2x3x4x5x6_share2_reg =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x6_share_in   ;
assign x0x1x2x3x4x5x7_share2_reg =  x0_share_in & x1_share_in & x2_share_in & x3_share_in & x4_share_in & x5_share_in & x7_share_in   ;



// second share of Degree-1 terms

assign x0_second_share = x0_subscript0_share2_reg ;
assign x1_second_share = x1_subscript0_share2_reg ;
assign x2_second_share = x2_subscript0_share2_reg ;
assign x3_second_share = x3_subscript0_share2_reg ;
assign x4_second_share = x4_subscript0_share2_reg ;
assign x5_second_share = x5_subscript0_share2_reg ;
assign x6_second_share = x6_subscript0_share2_reg ;
assign x7_second_share = x7_subscript0_share2_reg ;

// second share of Degree-2 terms

assign x0x1_second_share =  (x1_share2_reg  & x0_subscript0_share2_reg) ^ (x0_share2_reg  & x1_subscript0_share2_reg) ^ x0x1_subscript0_share2_reg ;
assign x0x2_second_share =  (x2_share2_reg  & x0_subscript0_share2_reg) ^ (x0_share2_reg  & x2_subscript0_share2_reg) ^ x0x2_subscript0_share2_reg ;
assign x0x3_second_share =  (x3_share2_reg  & x0_subscript0_share2_reg) ^ (x0_share2_reg  & x3_subscript0_share2_reg) ^ x0x3_subscript0_share2_reg ;
assign x0x4_second_share =  (x4_share2_reg  & x0_subscript0_share2_reg) ^ (x0_share2_reg  & x4_subscript0_share2_reg) ^ x0x4_subscript0_share2_reg ;
assign x0x5_second_share =  (x5_share2_reg  & x0_subscript0_share2_reg) ^ (x0_share2_reg  & x5_subscript0_share2_reg) ^ x0x5_subscript0_share2_reg ;
assign x0x6_second_share =  (x6_share2_reg  & x0_subscript0_share2_reg) ^ (x0_share2_reg  & x6_subscript0_share2_reg) ^ x0x6_subscript0_share2_reg ;
assign x0x7_second_share =  (x7_share2_reg  & x0_subscript0_share2_reg) ^ (x0_share2_reg  & x7_subscript0_share2_reg) ^ x0x7_subscript0_share2_reg ;
assign x1x2_second_share =  (x2_share2_reg  & x1_subscript0_share2_reg) ^ (x1_share2_reg  & x2_subscript0_share2_reg) ^ x1x2_subscript0_share2_reg ;
assign x1x3_second_share =  (x3_share2_reg  & x1_subscript0_share2_reg) ^ (x1_share2_reg  & x3_subscript0_share2_reg) ^ x1x3_subscript0_share2_reg ;
assign x1x4_second_share =  (x4_share2_reg  & x1_subscript0_share2_reg) ^ (x1_share2_reg  & x4_subscript0_share2_reg) ^ x1x4_subscript0_share2_reg ;
assign x1x5_second_share =  (x5_share2_reg  & x1_subscript0_share2_reg) ^ (x1_share2_reg  & x5_subscript0_share2_reg) ^ x1x5_subscript0_share2_reg ;
assign x1x6_second_share =  (x6_share2_reg  & x1_subscript0_share2_reg) ^ (x1_share2_reg  & x6_subscript0_share2_reg) ^ x1x6_subscript0_share2_reg ;
assign x1x7_second_share =  (x7_share2_reg  & x1_subscript0_share2_reg) ^ (x1_share2_reg  & x7_subscript0_share2_reg) ^ x1x7_subscript0_share2_reg ;
assign x2x3_second_share =  (x3_share2_reg  & x2_subscript0_share2_reg) ^ (x2_share2_reg  & x3_subscript0_share2_reg) ^ x2x3_subscript0_share2_reg ;
assign x2x4_second_share =  (x4_share2_reg  & x2_subscript0_share2_reg) ^ (x2_share2_reg  & x4_subscript0_share2_reg) ^ x2x4_subscript0_share2_reg ;
assign x2x5_second_share =  (x5_share2_reg  & x2_subscript0_share2_reg) ^ (x2_share2_reg  & x5_subscript0_share2_reg) ^ x2x5_subscript0_share2_reg ;
assign x2x6_second_share =  (x6_share2_reg  & x2_subscript0_share2_reg) ^ (x2_share2_reg  & x6_subscript0_share2_reg) ^ x2x6_subscript0_share2_reg ;
assign x2x7_second_share =  (x7_share2_reg  & x2_subscript0_share2_reg) ^ (x2_share2_reg  & x7_subscript0_share2_reg) ^ x2x7_subscript0_share2_reg ;
assign x3x4_second_share =  (x4_share2_reg  & x3_subscript0_share2_reg) ^ (x3_share2_reg  & x4_subscript0_share2_reg) ^ x3x4_subscript0_share2_reg ;
assign x3x5_second_share =  (x5_share2_reg  & x3_subscript0_share2_reg) ^ (x3_share2_reg  & x5_subscript0_share2_reg) ^ x3x5_subscript0_share2_reg ;
assign x3x6_second_share =  (x6_share2_reg  & x3_subscript0_share2_reg) ^ (x3_share2_reg  & x6_subscript0_share2_reg) ^ x3x6_subscript0_share2_reg ;
assign x3x7_second_share =  (x7_share2_reg  & x3_subscript0_share2_reg) ^ (x3_share2_reg  & x7_subscript0_share2_reg) ^ x3x7_subscript0_share2_reg ;
assign x4x5_second_share =  (x5_share2_reg  & x4_subscript0_share2_reg) ^ (x4_share2_reg  & x5_subscript0_share2_reg) ^ x4x5_subscript0_share2_reg ;
assign x4x6_second_share =  (x6_share2_reg  & x4_subscript0_share2_reg) ^ (x4_share2_reg  & x6_subscript0_share2_reg) ^ x4x6_subscript0_share2_reg ;
assign x4x7_second_share =  (x7_share2_reg  & x4_subscript0_share2_reg) ^ (x4_share2_reg  & x7_subscript0_share2_reg) ^ x4x7_subscript0_share2_reg ;
assign x5x6_second_share =  (x6_share2_reg  & x5_subscript0_share2_reg) ^ (x5_share2_reg  & x6_subscript0_share2_reg) ^ x5x6_subscript0_share2_reg ;
assign x5x7_second_share =  (x7_share2_reg  & x5_subscript0_share2_reg) ^ (x5_share2_reg  & x7_subscript0_share2_reg) ^ x5x7_subscript0_share2_reg ;
assign x6x7_second_share =  (x7_share2_reg  & x6_subscript0_share2_reg) ^ (x6_share2_reg  & x7_subscript0_share2_reg) ^ x6x7_subscript0_share2_reg ;


// second share of Degree-3 terms

assign x0x1x2_second_share =  x0_share2_reg & x1x2_second_share ^x1x2_share2_reg  & x0_subscript0_share2_reg ^ x2_share2_reg  & x0x1_subscript0_share2_reg ^ x1_share2_reg  & x0x2_subscript0_share2_reg ^ x0x1x2_subscript0_share2_reg ;
assign x0x1x3_second_share =  x0_share2_reg & x1x3_second_share ^x1x3_share2_reg  & x0_subscript0_share2_reg ^ x3_share2_reg  & x0x1_subscript0_share2_reg ^ x1_share2_reg  & x0x3_subscript0_share2_reg ^ x0x1x3_subscript0_share2_reg ;
assign x0x1x4_second_share =  x0_share2_reg & x1x4_second_share ^x1x4_share2_reg  & x0_subscript0_share2_reg ^ x4_share2_reg  & x0x1_subscript0_share2_reg ^ x1_share2_reg  & x0x4_subscript0_share2_reg ^ x0x1x4_subscript0_share2_reg ;
assign x0x1x5_second_share =  x0_share2_reg & x1x5_second_share ^x1x5_share2_reg  & x0_subscript0_share2_reg ^ x5_share2_reg  & x0x1_subscript0_share2_reg ^ x1_share2_reg  & x0x5_subscript0_share2_reg ^ x0x1x5_subscript0_share2_reg ;
assign x0x1x6_second_share =  x0_share2_reg & x1x6_second_share ^x1x6_share2_reg  & x0_subscript0_share2_reg ^ x6_share2_reg  & x0x1_subscript0_share2_reg ^ x1_share2_reg  & x0x6_subscript0_share2_reg ^ x0x1x6_subscript0_share2_reg ;
assign x0x1x7_second_share =  x0_share2_reg & x1x7_second_share ^x1x7_share2_reg  & x0_subscript0_share2_reg ^ x7_share2_reg  & x0x1_subscript0_share2_reg ^ x1_share2_reg  & x0x7_subscript0_share2_reg ^ x0x1x7_subscript0_share2_reg ;
assign x0x2x3_second_share =  x0_share2_reg & x2x3_second_share ^x2x3_share2_reg  & x0_subscript0_share2_reg ^ x3_share2_reg  & x0x2_subscript0_share2_reg ^ x2_share2_reg  & x0x3_subscript0_share2_reg ^ x0x2x3_subscript0_share2_reg ;
assign x0x2x4_second_share =  x0_share2_reg & x2x4_second_share ^x2x4_share2_reg  & x0_subscript0_share2_reg ^ x4_share2_reg  & x0x2_subscript0_share2_reg ^ x2_share2_reg  & x0x4_subscript0_share2_reg ^ x0x2x4_subscript0_share2_reg ;
assign x0x2x5_second_share =  x0_share2_reg & x2x5_second_share ^x2x5_share2_reg  & x0_subscript0_share2_reg ^ x5_share2_reg  & x0x2_subscript0_share2_reg ^ x2_share2_reg  & x0x5_subscript0_share2_reg ^ x0x2x5_subscript0_share2_reg ;
assign x0x2x6_second_share =  x0_share2_reg & x2x6_second_share ^x2x6_share2_reg  & x0_subscript0_share2_reg ^ x6_share2_reg  & x0x2_subscript0_share2_reg ^ x2_share2_reg  & x0x6_subscript0_share2_reg ^ x0x2x6_subscript0_share2_reg ;
assign x0x2x7_second_share =  x0_share2_reg & x2x7_second_share ^x2x7_share2_reg  & x0_subscript0_share2_reg ^ x7_share2_reg  & x0x2_subscript0_share2_reg ^ x2_share2_reg  & x0x7_subscript0_share2_reg ^ x0x2x7_subscript0_share2_reg ;
assign x0x3x4_second_share =  x0_share2_reg & x3x4_second_share ^x3x4_share2_reg  & x0_subscript0_share2_reg ^ x4_share2_reg  & x0x3_subscript0_share2_reg ^ x3_share2_reg  & x0x4_subscript0_share2_reg ^ x0x3x4_subscript0_share2_reg ;
assign x0x3x5_second_share =  x0_share2_reg & x3x5_second_share ^x3x5_share2_reg  & x0_subscript0_share2_reg ^ x5_share2_reg  & x0x3_subscript0_share2_reg ^ x3_share2_reg  & x0x5_subscript0_share2_reg ^ x0x3x5_subscript0_share2_reg ;
assign x0x3x6_second_share =  x0_share2_reg & x3x6_second_share ^x3x6_share2_reg  & x0_subscript0_share2_reg ^ x6_share2_reg  & x0x3_subscript0_share2_reg ^ x3_share2_reg  & x0x6_subscript0_share2_reg ^ x0x3x6_subscript0_share2_reg ;
assign x0x3x7_second_share =  x0_share2_reg & x3x7_second_share ^x3x7_share2_reg  & x0_subscript0_share2_reg ^ x7_share2_reg  & x0x3_subscript0_share2_reg ^ x3_share2_reg  & x0x7_subscript0_share2_reg ^ x0x3x7_subscript0_share2_reg ;
assign x0x4x5_second_share =  x0_share2_reg & x4x5_second_share ^x4x5_share2_reg  & x0_subscript0_share2_reg ^ x5_share2_reg  & x0x4_subscript0_share2_reg ^ x4_share2_reg  & x0x5_subscript0_share2_reg ^ x0x4x5_subscript0_share2_reg ;
assign x0x4x6_second_share =  x0_share2_reg & x4x6_second_share ^x4x6_share2_reg  & x0_subscript0_share2_reg ^ x6_share2_reg  & x0x4_subscript0_share2_reg ^ x4_share2_reg  & x0x6_subscript0_share2_reg ^ x0x4x6_subscript0_share2_reg ;
assign x0x4x7_second_share =  x0_share2_reg & x4x7_second_share ^x4x7_share2_reg  & x0_subscript0_share2_reg ^ x7_share2_reg  & x0x4_subscript0_share2_reg ^ x4_share2_reg  & x0x7_subscript0_share2_reg ^ x0x4x7_subscript0_share2_reg ;
assign x0x5x6_second_share =  x0_share2_reg & x5x6_second_share ^x5x6_share2_reg  & x0_subscript0_share2_reg ^ x6_share2_reg  & x0x5_subscript0_share2_reg ^ x5_share2_reg  & x0x6_subscript0_share2_reg ^ x0x5x6_subscript0_share2_reg ;
assign x0x5x7_second_share =  x0_share2_reg & x5x7_second_share ^x5x7_share2_reg  & x0_subscript0_share2_reg ^ x7_share2_reg  & x0x5_subscript0_share2_reg ^ x5_share2_reg  & x0x7_subscript0_share2_reg ^ x0x5x7_subscript0_share2_reg ;
assign x0x6x7_second_share =  x0_share2_reg & x6x7_second_share ^x6x7_share2_reg  & x0_subscript0_share2_reg ^ x7_share2_reg  & x0x6_subscript0_share2_reg ^ x6_share2_reg  & x0x7_subscript0_share2_reg ^ x0x6x7_subscript0_share2_reg ;
assign x1x2x3_second_share =  x1_share2_reg & x2x3_second_share ^x2x3_share2_reg  & x1_subscript0_share2_reg ^ x3_share2_reg  & x1x2_subscript0_share2_reg ^ x2_share2_reg  & x1x3_subscript0_share2_reg ^ x1x2x3_subscript0_share2_reg ;
assign x1x2x4_second_share =  x1_share2_reg & x2x4_second_share ^x2x4_share2_reg  & x1_subscript0_share2_reg ^ x4_share2_reg  & x1x2_subscript0_share2_reg ^ x2_share2_reg  & x1x4_subscript0_share2_reg ^ x1x2x4_subscript0_share2_reg ;
assign x1x2x5_second_share =  x1_share2_reg & x2x5_second_share ^x2x5_share2_reg  & x1_subscript0_share2_reg ^ x5_share2_reg  & x1x2_subscript0_share2_reg ^ x2_share2_reg  & x1x5_subscript0_share2_reg ^ x1x2x5_subscript0_share2_reg ;
assign x1x2x6_second_share =  x1_share2_reg & x2x6_second_share ^x2x6_share2_reg  & x1_subscript0_share2_reg ^ x6_share2_reg  & x1x2_subscript0_share2_reg ^ x2_share2_reg  & x1x6_subscript0_share2_reg ^ x1x2x6_subscript0_share2_reg ;
assign x1x2x7_second_share =  x1_share2_reg & x2x7_second_share ^x2x7_share2_reg  & x1_subscript0_share2_reg ^ x7_share2_reg  & x1x2_subscript0_share2_reg ^ x2_share2_reg  & x1x7_subscript0_share2_reg ^ x1x2x7_subscript0_share2_reg ;
assign x1x3x4_second_share =  x1_share2_reg & x3x4_second_share ^x3x4_share2_reg  & x1_subscript0_share2_reg ^ x4_share2_reg  & x1x3_subscript0_share2_reg ^ x3_share2_reg  & x1x4_subscript0_share2_reg ^ x1x3x4_subscript0_share2_reg ;
assign x1x3x5_second_share =  x1_share2_reg & x3x5_second_share ^x3x5_share2_reg  & x1_subscript0_share2_reg ^ x5_share2_reg  & x1x3_subscript0_share2_reg ^ x3_share2_reg  & x1x5_subscript0_share2_reg ^ x1x3x5_subscript0_share2_reg ;
assign x1x3x6_second_share =  x1_share2_reg & x3x6_second_share ^x3x6_share2_reg  & x1_subscript0_share2_reg ^ x6_share2_reg  & x1x3_subscript0_share2_reg ^ x3_share2_reg  & x1x6_subscript0_share2_reg ^ x1x3x6_subscript0_share2_reg ;
assign x1x3x7_second_share =  x1_share2_reg & x3x7_second_share ^x3x7_share2_reg  & x1_subscript0_share2_reg ^ x7_share2_reg  & x1x3_subscript0_share2_reg ^ x3_share2_reg  & x1x7_subscript0_share2_reg ^ x1x3x7_subscript0_share2_reg ;
assign x1x4x5_second_share =  x1_share2_reg & x4x5_second_share ^x4x5_share2_reg  & x1_subscript0_share2_reg ^ x5_share2_reg  & x1x4_subscript0_share2_reg ^ x4_share2_reg  & x1x5_subscript0_share2_reg ^ x1x4x5_subscript0_share2_reg ;
assign x1x4x6_second_share =  x1_share2_reg & x4x6_second_share ^x4x6_share2_reg  & x1_subscript0_share2_reg ^ x6_share2_reg  & x1x4_subscript0_share2_reg ^ x4_share2_reg  & x1x6_subscript0_share2_reg ^ x1x4x6_subscript0_share2_reg ;
assign x1x4x7_second_share =  x1_share2_reg & x4x7_second_share ^x4x7_share2_reg  & x1_subscript0_share2_reg ^ x7_share2_reg  & x1x4_subscript0_share2_reg ^ x4_share2_reg  & x1x7_subscript0_share2_reg ^ x1x4x7_subscript0_share2_reg ;
assign x1x5x6_second_share =  x1_share2_reg & x5x6_second_share ^x5x6_share2_reg  & x1_subscript0_share2_reg ^ x6_share2_reg  & x1x5_subscript0_share2_reg ^ x5_share2_reg  & x1x6_subscript0_share2_reg ^ x1x5x6_subscript0_share2_reg ;
assign x1x5x7_second_share =  x1_share2_reg & x5x7_second_share ^x5x7_share2_reg  & x1_subscript0_share2_reg ^ x7_share2_reg  & x1x5_subscript0_share2_reg ^ x5_share2_reg  & x1x7_subscript0_share2_reg ^ x1x5x7_subscript0_share2_reg ;
assign x1x6x7_second_share =  x1_share2_reg & x6x7_second_share ^x6x7_share2_reg  & x1_subscript0_share2_reg ^ x7_share2_reg  & x1x6_subscript0_share2_reg ^ x6_share2_reg  & x1x7_subscript0_share2_reg ^ x1x6x7_subscript0_share2_reg ;
assign x2x3x4_second_share =  x2_share2_reg & x3x4_second_share ^x3x4_share2_reg  & x2_subscript0_share2_reg ^ x4_share2_reg  & x2x3_subscript0_share2_reg ^ x3_share2_reg  & x2x4_subscript0_share2_reg ^ x2x3x4_subscript0_share2_reg ;
assign x2x3x5_second_share =  x2_share2_reg & x3x5_second_share ^x3x5_share2_reg  & x2_subscript0_share2_reg ^ x5_share2_reg  & x2x3_subscript0_share2_reg ^ x3_share2_reg  & x2x5_subscript0_share2_reg ^ x2x3x5_subscript0_share2_reg ;
assign x2x3x6_second_share =  x2_share2_reg & x3x6_second_share ^x3x6_share2_reg  & x2_subscript0_share2_reg ^ x6_share2_reg  & x2x3_subscript0_share2_reg ^ x3_share2_reg  & x2x6_subscript0_share2_reg ^ x2x3x6_subscript0_share2_reg ;
assign x2x3x7_second_share =  x2_share2_reg & x3x7_second_share ^x3x7_share2_reg  & x2_subscript0_share2_reg ^ x7_share2_reg  & x2x3_subscript0_share2_reg ^ x3_share2_reg  & x2x7_subscript0_share2_reg ^ x2x3x7_subscript0_share2_reg ;
assign x2x4x5_second_share =  x2_share2_reg & x4x5_second_share ^x4x5_share2_reg  & x2_subscript0_share2_reg ^ x5_share2_reg  & x2x4_subscript0_share2_reg ^ x4_share2_reg  & x2x5_subscript0_share2_reg ^ x2x4x5_subscript0_share2_reg ;
assign x2x4x6_second_share =  x2_share2_reg & x4x6_second_share ^x4x6_share2_reg  & x2_subscript0_share2_reg ^ x6_share2_reg  & x2x4_subscript0_share2_reg ^ x4_share2_reg  & x2x6_subscript0_share2_reg ^ x2x4x6_subscript0_share2_reg ;
assign x2x4x7_second_share =  x2_share2_reg & x4x7_second_share ^x4x7_share2_reg  & x2_subscript0_share2_reg ^ x7_share2_reg  & x2x4_subscript0_share2_reg ^ x4_share2_reg  & x2x7_subscript0_share2_reg ^ x2x4x7_subscript0_share2_reg ;
assign x2x5x6_second_share =  x2_share2_reg & x5x6_second_share ^x5x6_share2_reg  & x2_subscript0_share2_reg ^ x6_share2_reg  & x2x5_subscript0_share2_reg ^ x5_share2_reg  & x2x6_subscript0_share2_reg ^ x2x5x6_subscript0_share2_reg ;
assign x2x5x7_second_share =  x2_share2_reg & x5x7_second_share ^x5x7_share2_reg  & x2_subscript0_share2_reg ^ x7_share2_reg  & x2x5_subscript0_share2_reg ^ x5_share2_reg  & x2x7_subscript0_share2_reg ^ x2x5x7_subscript0_share2_reg ;
assign x2x6x7_second_share =  x2_share2_reg & x6x7_second_share ^x6x7_share2_reg  & x2_subscript0_share2_reg ^ x7_share2_reg  & x2x6_subscript0_share2_reg ^ x6_share2_reg  & x2x7_subscript0_share2_reg ^ x2x6x7_subscript0_share2_reg ;
assign x3x4x5_second_share =  x3_share2_reg & x4x5_second_share ^x4x5_share2_reg  & x3_subscript0_share2_reg ^ x5_share2_reg  & x3x4_subscript0_share2_reg ^ x4_share2_reg  & x3x5_subscript0_share2_reg ^ x3x4x5_subscript0_share2_reg ;
assign x3x4x6_second_share =  x3_share2_reg & x4x6_second_share ^x4x6_share2_reg  & x3_subscript0_share2_reg ^ x6_share2_reg  & x3x4_subscript0_share2_reg ^ x4_share2_reg  & x3x6_subscript0_share2_reg ^ x3x4x6_subscript0_share2_reg ;
assign x3x4x7_second_share =  x3_share2_reg & x4x7_second_share ^x4x7_share2_reg  & x3_subscript0_share2_reg ^ x7_share2_reg  & x3x4_subscript0_share2_reg ^ x4_share2_reg  & x3x7_subscript0_share2_reg ^ x3x4x7_subscript0_share2_reg ;
assign x3x5x6_second_share =  x3_share2_reg & x5x6_second_share ^x5x6_share2_reg  & x3_subscript0_share2_reg ^ x6_share2_reg  & x3x5_subscript0_share2_reg ^ x5_share2_reg  & x3x6_subscript0_share2_reg ^ x3x5x6_subscript0_share2_reg ;
assign x3x5x7_second_share =  x3_share2_reg & x5x7_second_share ^x5x7_share2_reg  & x3_subscript0_share2_reg ^ x7_share2_reg  & x3x5_subscript0_share2_reg ^ x5_share2_reg  & x3x7_subscript0_share2_reg ^ x3x5x7_subscript0_share2_reg ;
assign x3x6x7_second_share =  x3_share2_reg & x6x7_second_share ^x6x7_share2_reg  & x3_subscript0_share2_reg ^ x7_share2_reg  & x3x6_subscript0_share2_reg ^ x6_share2_reg  & x3x7_subscript0_share2_reg ^ x3x6x7_subscript0_share2_reg ;
assign x4x5x6_second_share =  x4_share2_reg & x5x6_second_share ^x5x6_share2_reg  & x4_subscript0_share2_reg ^ x6_share2_reg  & x4x5_subscript0_share2_reg ^ x5_share2_reg  & x4x6_subscript0_share2_reg ^ x4x5x6_subscript0_share2_reg ;
assign x4x5x7_second_share =  x4_share2_reg & x5x7_second_share ^x5x7_share2_reg  & x4_subscript0_share2_reg ^ x7_share2_reg  & x4x5_subscript0_share2_reg ^ x5_share2_reg  & x4x7_subscript0_share2_reg ^ x4x5x7_subscript0_share2_reg ;
assign x4x6x7_second_share =  x4_share2_reg & x6x7_second_share ^x6x7_share2_reg  & x4_subscript0_share2_reg ^ x7_share2_reg  & x4x6_subscript0_share2_reg ^ x6_share2_reg  & x4x7_subscript0_share2_reg ^ x4x6x7_subscript0_share2_reg ;
assign x5x6x7_second_share =  x5_share2_reg & x6x7_second_share ^x6x7_share2_reg  & x5_subscript0_share2_reg ^ x7_share2_reg  & x5x6_subscript0_share2_reg ^ x6_share2_reg  & x5x7_subscript0_share2_reg ^ x5x6x7_subscript0_share2_reg ;


// second share of Degree-4 terms


assign x0x1x2x3_second_share =      x0_share2_reg & x1x2x3_second_share ^    x1_share2_reg & x0x2x3_second_share ^    x0x1_share2_reg  & x2x3_second_share ^     x2_share2_reg  & x0x1x3_subscript0_share2_reg ^ x3_share2_reg  & x0x1x2_subscript0_share2_reg ^    x2x3_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x2x3_subscript0_share2_reg ;
assign x0x1x2x4_second_share =      x0_share2_reg & x1x2x4_second_share ^    x1_share2_reg & x0x2x4_second_share ^    x0x1_share2_reg  & x2x4_second_share ^     x2_share2_reg  & x0x1x4_subscript0_share2_reg ^ x4_share2_reg  & x0x1x2_subscript0_share2_reg ^    x2x4_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x2x4_subscript0_share2_reg ;
assign x0x1x2x5_second_share =      x0_share2_reg & x1x2x5_second_share ^    x1_share2_reg & x0x2x5_second_share ^    x0x1_share2_reg  & x2x5_second_share ^     x2_share2_reg  & x0x1x5_subscript0_share2_reg ^ x5_share2_reg  & x0x1x2_subscript0_share2_reg ^    x2x5_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x2x5_subscript0_share2_reg ;
assign x0x1x2x6_second_share =      x0_share2_reg & x1x2x6_second_share ^    x1_share2_reg & x0x2x6_second_share ^    x0x1_share2_reg  & x2x6_second_share ^     x2_share2_reg  & x0x1x6_subscript0_share2_reg ^ x6_share2_reg  & x0x1x2_subscript0_share2_reg ^    x2x6_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x2x6_subscript0_share2_reg ;
assign x0x1x2x7_second_share =      x0_share2_reg & x1x2x7_second_share ^    x1_share2_reg & x0x2x7_second_share ^    x0x1_share2_reg  & x2x7_second_share ^     x2_share2_reg  & x0x1x7_subscript0_share2_reg ^ x7_share2_reg  & x0x1x2_subscript0_share2_reg ^    x2x7_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x2x7_subscript0_share2_reg ;
assign x0x1x3x4_second_share =      x0_share2_reg & x1x3x4_second_share ^    x1_share2_reg & x0x3x4_second_share ^    x0x1_share2_reg  & x3x4_second_share ^     x3_share2_reg  & x0x1x4_subscript0_share2_reg ^ x4_share2_reg  & x0x1x3_subscript0_share2_reg ^    x3x4_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x3x4_subscript0_share2_reg ;
assign x0x1x3x5_second_share =      x0_share2_reg & x1x3x5_second_share ^    x1_share2_reg & x0x3x5_second_share ^    x0x1_share2_reg  & x3x5_second_share ^     x3_share2_reg  & x0x1x5_subscript0_share2_reg ^ x5_share2_reg  & x0x1x3_subscript0_share2_reg ^    x3x5_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x3x5_subscript0_share2_reg ;
assign x0x1x3x6_second_share =      x0_share2_reg & x1x3x6_second_share ^    x1_share2_reg & x0x3x6_second_share ^    x0x1_share2_reg  & x3x6_second_share ^     x3_share2_reg  & x0x1x6_subscript0_share2_reg ^ x6_share2_reg  & x0x1x3_subscript0_share2_reg ^    x3x6_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x3x6_subscript0_share2_reg ;
assign x0x1x3x7_second_share =      x0_share2_reg & x1x3x7_second_share ^    x1_share2_reg & x0x3x7_second_share ^    x0x1_share2_reg  & x3x7_second_share ^     x3_share2_reg  & x0x1x7_subscript0_share2_reg ^ x7_share2_reg  & x0x1x3_subscript0_share2_reg ^    x3x7_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x3x7_subscript0_share2_reg ;
assign x0x1x4x5_second_share =      x0_share2_reg & x1x4x5_second_share ^    x1_share2_reg & x0x4x5_second_share ^    x0x1_share2_reg  & x4x5_second_share ^     x4_share2_reg  & x0x1x5_subscript0_share2_reg ^ x5_share2_reg  & x0x1x4_subscript0_share2_reg ^    x4x5_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x4x5_subscript0_share2_reg ;
assign x0x1x4x6_second_share =      x0_share2_reg & x1x4x6_second_share ^    x1_share2_reg & x0x4x6_second_share ^    x0x1_share2_reg  & x4x6_second_share ^     x4_share2_reg  & x0x1x6_subscript0_share2_reg ^ x6_share2_reg  & x0x1x4_subscript0_share2_reg ^    x4x6_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x4x6_subscript0_share2_reg ;
assign x0x1x4x7_second_share =      x0_share2_reg & x1x4x7_second_share ^    x1_share2_reg & x0x4x7_second_share ^    x0x1_share2_reg  & x4x7_second_share ^     x4_share2_reg  & x0x1x7_subscript0_share2_reg ^ x7_share2_reg  & x0x1x4_subscript0_share2_reg ^    x4x7_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x4x7_subscript0_share2_reg ;
assign x0x1x5x6_second_share =      x0_share2_reg & x1x5x6_second_share ^    x1_share2_reg & x0x5x6_second_share ^    x0x1_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x0x1x6_subscript0_share2_reg ^ x6_share2_reg  & x0x1x5_subscript0_share2_reg ^    x5x6_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x5x6_subscript0_share2_reg ;
assign x0x1x5x7_second_share =      x0_share2_reg & x1x5x7_second_share ^    x1_share2_reg & x0x5x7_second_share ^    x0x1_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x0x1x7_subscript0_share2_reg ^ x7_share2_reg  & x0x1x5_subscript0_share2_reg ^    x5x7_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x5x7_subscript0_share2_reg ;
assign x0x1x6x7_second_share =      x0_share2_reg & x1x6x7_second_share ^    x1_share2_reg & x0x6x7_second_share ^    x0x1_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x0x1x7_subscript0_share2_reg ^ x7_share2_reg  & x0x1x6_subscript0_share2_reg ^    x6x7_share2_reg  & x0x1_subscript0_share2_reg ^x0x1x6x7_subscript0_share2_reg ;
assign x0x2x3x4_second_share =      x0_share2_reg & x2x3x4_second_share ^    x2_share2_reg & x0x3x4_second_share ^    x0x2_share2_reg  & x3x4_second_share ^     x3_share2_reg  & x0x2x4_subscript0_share2_reg ^ x4_share2_reg  & x0x2x3_subscript0_share2_reg ^    x3x4_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x3x4_subscript0_share2_reg ;
assign x0x2x3x5_second_share =      x0_share2_reg & x2x3x5_second_share ^    x2_share2_reg & x0x3x5_second_share ^    x0x2_share2_reg  & x3x5_second_share ^     x3_share2_reg  & x0x2x5_subscript0_share2_reg ^ x5_share2_reg  & x0x2x3_subscript0_share2_reg ^    x3x5_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x3x5_subscript0_share2_reg ;
assign x0x2x3x6_second_share =      x0_share2_reg & x2x3x6_second_share ^    x2_share2_reg & x0x3x6_second_share ^    x0x2_share2_reg  & x3x6_second_share ^     x3_share2_reg  & x0x2x6_subscript0_share2_reg ^ x6_share2_reg  & x0x2x3_subscript0_share2_reg ^    x3x6_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x3x6_subscript0_share2_reg ;
assign x0x2x3x7_second_share =      x0_share2_reg & x2x3x7_second_share ^    x2_share2_reg & x0x3x7_second_share ^    x0x2_share2_reg  & x3x7_second_share ^     x3_share2_reg  & x0x2x7_subscript0_share2_reg ^ x7_share2_reg  & x0x2x3_subscript0_share2_reg ^    x3x7_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x3x7_subscript0_share2_reg ;
assign x0x2x4x5_second_share =      x0_share2_reg & x2x4x5_second_share ^    x2_share2_reg & x0x4x5_second_share ^    x0x2_share2_reg  & x4x5_second_share ^     x4_share2_reg  & x0x2x5_subscript0_share2_reg ^ x5_share2_reg  & x0x2x4_subscript0_share2_reg ^    x4x5_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x4x5_subscript0_share2_reg ;
assign x0x2x4x6_second_share =      x0_share2_reg & x2x4x6_second_share ^    x2_share2_reg & x0x4x6_second_share ^    x0x2_share2_reg  & x4x6_second_share ^     x4_share2_reg  & x0x2x6_subscript0_share2_reg ^ x6_share2_reg  & x0x2x4_subscript0_share2_reg ^    x4x6_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x4x6_subscript0_share2_reg ;
assign x0x2x4x7_second_share =      x0_share2_reg & x2x4x7_second_share ^    x2_share2_reg & x0x4x7_second_share ^    x0x2_share2_reg  & x4x7_second_share ^     x4_share2_reg  & x0x2x7_subscript0_share2_reg ^ x7_share2_reg  & x0x2x4_subscript0_share2_reg ^    x4x7_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x4x7_subscript0_share2_reg ;
assign x0x2x5x6_second_share =      x0_share2_reg & x2x5x6_second_share ^    x2_share2_reg & x0x5x6_second_share ^    x0x2_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x0x2x6_subscript0_share2_reg ^ x6_share2_reg  & x0x2x5_subscript0_share2_reg ^    x5x6_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x5x6_subscript0_share2_reg ;
assign x0x2x5x7_second_share =      x0_share2_reg & x2x5x7_second_share ^    x2_share2_reg & x0x5x7_second_share ^    x0x2_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x0x2x7_subscript0_share2_reg ^ x7_share2_reg  & x0x2x5_subscript0_share2_reg ^    x5x7_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x5x7_subscript0_share2_reg ;
assign x0x2x6x7_second_share =      x0_share2_reg & x2x6x7_second_share ^    x2_share2_reg & x0x6x7_second_share ^    x0x2_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x0x2x7_subscript0_share2_reg ^ x7_share2_reg  & x0x2x6_subscript0_share2_reg ^    x6x7_share2_reg  & x0x2_subscript0_share2_reg ^x0x2x6x7_subscript0_share2_reg ;
assign x0x3x4x5_second_share =      x0_share2_reg & x3x4x5_second_share ^    x3_share2_reg & x0x4x5_second_share ^    x0x3_share2_reg  & x4x5_second_share ^     x4_share2_reg  & x0x3x5_subscript0_share2_reg ^ x5_share2_reg  & x0x3x4_subscript0_share2_reg ^    x4x5_share2_reg  & x0x3_subscript0_share2_reg ^x0x3x4x5_subscript0_share2_reg ;
assign x0x3x4x6_second_share =      x0_share2_reg & x3x4x6_second_share ^    x3_share2_reg & x0x4x6_second_share ^    x0x3_share2_reg  & x4x6_second_share ^     x4_share2_reg  & x0x3x6_subscript0_share2_reg ^ x6_share2_reg  & x0x3x4_subscript0_share2_reg ^    x4x6_share2_reg  & x0x3_subscript0_share2_reg ^x0x3x4x6_subscript0_share2_reg ;
assign x0x3x4x7_second_share =      x0_share2_reg & x3x4x7_second_share ^    x3_share2_reg & x0x4x7_second_share ^    x0x3_share2_reg  & x4x7_second_share ^     x4_share2_reg  & x0x3x7_subscript0_share2_reg ^ x7_share2_reg  & x0x3x4_subscript0_share2_reg ^    x4x7_share2_reg  & x0x3_subscript0_share2_reg ^x0x3x4x7_subscript0_share2_reg ;
assign x0x3x5x6_second_share =      x0_share2_reg & x3x5x6_second_share ^    x3_share2_reg & x0x5x6_second_share ^    x0x3_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x0x3x6_subscript0_share2_reg ^ x6_share2_reg  & x0x3x5_subscript0_share2_reg ^    x5x6_share2_reg  & x0x3_subscript0_share2_reg ^x0x3x5x6_subscript0_share2_reg ;
assign x0x3x5x7_second_share =      x0_share2_reg & x3x5x7_second_share ^    x3_share2_reg & x0x5x7_second_share ^    x0x3_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x0x3x7_subscript0_share2_reg ^ x7_share2_reg  & x0x3x5_subscript0_share2_reg ^    x5x7_share2_reg  & x0x3_subscript0_share2_reg ^x0x3x5x7_subscript0_share2_reg ;
assign x0x3x6x7_second_share =      x0_share2_reg & x3x6x7_second_share ^    x3_share2_reg & x0x6x7_second_share ^    x0x3_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x0x3x7_subscript0_share2_reg ^ x7_share2_reg  & x0x3x6_subscript0_share2_reg ^    x6x7_share2_reg  & x0x3_subscript0_share2_reg ^x0x3x6x7_subscript0_share2_reg ;
assign x0x4x5x6_second_share =      x0_share2_reg & x4x5x6_second_share ^    x4_share2_reg & x0x5x6_second_share ^    x0x4_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x0x4x6_subscript0_share2_reg ^ x6_share2_reg  & x0x4x5_subscript0_share2_reg ^    x5x6_share2_reg  & x0x4_subscript0_share2_reg ^x0x4x5x6_subscript0_share2_reg ;
assign x0x4x5x7_second_share =      x0_share2_reg & x4x5x7_second_share ^    x4_share2_reg & x0x5x7_second_share ^    x0x4_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x0x4x7_subscript0_share2_reg ^ x7_share2_reg  & x0x4x5_subscript0_share2_reg ^    x5x7_share2_reg  & x0x4_subscript0_share2_reg ^x0x4x5x7_subscript0_share2_reg ;
assign x0x4x6x7_second_share =      x0_share2_reg & x4x6x7_second_share ^    x4_share2_reg & x0x6x7_second_share ^    x0x4_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x0x4x7_subscript0_share2_reg ^ x7_share2_reg  & x0x4x6_subscript0_share2_reg ^    x6x7_share2_reg  & x0x4_subscript0_share2_reg ^x0x4x6x7_subscript0_share2_reg ;
assign x0x5x6x7_second_share =      x0_share2_reg & x5x6x7_second_share ^    x5_share2_reg & x0x6x7_second_share ^    x0x5_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x0x5x7_subscript0_share2_reg ^ x7_share2_reg  & x0x5x6_subscript0_share2_reg ^    x6x7_share2_reg  & x0x5_subscript0_share2_reg ^x0x5x6x7_subscript0_share2_reg ;
assign x1x2x3x4_second_share =      x1_share2_reg & x2x3x4_second_share ^    x2_share2_reg & x1x3x4_second_share ^    x1x2_share2_reg  & x3x4_second_share ^     x3_share2_reg  & x1x2x4_subscript0_share2_reg ^ x4_share2_reg  & x1x2x3_subscript0_share2_reg ^    x3x4_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x3x4_subscript0_share2_reg ;
assign x1x2x3x5_second_share =      x1_share2_reg & x2x3x5_second_share ^    x2_share2_reg & x1x3x5_second_share ^    x1x2_share2_reg  & x3x5_second_share ^     x3_share2_reg  & x1x2x5_subscript0_share2_reg ^ x5_share2_reg  & x1x2x3_subscript0_share2_reg ^    x3x5_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x3x5_subscript0_share2_reg ;
assign x1x2x3x6_second_share =      x1_share2_reg & x2x3x6_second_share ^    x2_share2_reg & x1x3x6_second_share ^    x1x2_share2_reg  & x3x6_second_share ^     x3_share2_reg  & x1x2x6_subscript0_share2_reg ^ x6_share2_reg  & x1x2x3_subscript0_share2_reg ^    x3x6_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x3x6_subscript0_share2_reg ;
assign x1x2x3x7_second_share =      x1_share2_reg & x2x3x7_second_share ^    x2_share2_reg & x1x3x7_second_share ^    x1x2_share2_reg  & x3x7_second_share ^     x3_share2_reg  & x1x2x7_subscript0_share2_reg ^ x7_share2_reg  & x1x2x3_subscript0_share2_reg ^    x3x7_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x3x7_subscript0_share2_reg ;
assign x1x2x4x5_second_share =      x1_share2_reg & x2x4x5_second_share ^    x2_share2_reg & x1x4x5_second_share ^    x1x2_share2_reg  & x4x5_second_share ^     x4_share2_reg  & x1x2x5_subscript0_share2_reg ^ x5_share2_reg  & x1x2x4_subscript0_share2_reg ^    x4x5_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x4x5_subscript0_share2_reg ;
assign x1x2x4x6_second_share =      x1_share2_reg & x2x4x6_second_share ^    x2_share2_reg & x1x4x6_second_share ^    x1x2_share2_reg  & x4x6_second_share ^     x4_share2_reg  & x1x2x6_subscript0_share2_reg ^ x6_share2_reg  & x1x2x4_subscript0_share2_reg ^    x4x6_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x4x6_subscript0_share2_reg ;
assign x1x2x4x7_second_share =      x1_share2_reg & x2x4x7_second_share ^    x2_share2_reg & x1x4x7_second_share ^    x1x2_share2_reg  & x4x7_second_share ^     x4_share2_reg  & x1x2x7_subscript0_share2_reg ^ x7_share2_reg  & x1x2x4_subscript0_share2_reg ^    x4x7_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x4x7_subscript0_share2_reg ;
assign x1x2x5x6_second_share =      x1_share2_reg & x2x5x6_second_share ^    x2_share2_reg & x1x5x6_second_share ^    x1x2_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x1x2x6_subscript0_share2_reg ^ x6_share2_reg  & x1x2x5_subscript0_share2_reg ^    x5x6_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x5x6_subscript0_share2_reg ;
assign x1x2x5x7_second_share =      x1_share2_reg & x2x5x7_second_share ^    x2_share2_reg & x1x5x7_second_share ^    x1x2_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x1x2x7_subscript0_share2_reg ^ x7_share2_reg  & x1x2x5_subscript0_share2_reg ^    x5x7_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x5x7_subscript0_share2_reg ;
assign x1x2x6x7_second_share =      x1_share2_reg & x2x6x7_second_share ^    x2_share2_reg & x1x6x7_second_share ^    x1x2_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x1x2x7_subscript0_share2_reg ^ x7_share2_reg  & x1x2x6_subscript0_share2_reg ^    x6x7_share2_reg  & x1x2_subscript0_share2_reg ^x1x2x6x7_subscript0_share2_reg ;
assign x1x3x4x5_second_share =      x1_share2_reg & x3x4x5_second_share ^    x3_share2_reg & x1x4x5_second_share ^    x1x3_share2_reg  & x4x5_second_share ^     x4_share2_reg  & x1x3x5_subscript0_share2_reg ^ x5_share2_reg  & x1x3x4_subscript0_share2_reg ^    x4x5_share2_reg  & x1x3_subscript0_share2_reg ^x1x3x4x5_subscript0_share2_reg ;
assign x1x3x4x6_second_share =      x1_share2_reg & x3x4x6_second_share ^    x3_share2_reg & x1x4x6_second_share ^    x1x3_share2_reg  & x4x6_second_share ^     x4_share2_reg  & x1x3x6_subscript0_share2_reg ^ x6_share2_reg  & x1x3x4_subscript0_share2_reg ^    x4x6_share2_reg  & x1x3_subscript0_share2_reg ^x1x3x4x6_subscript0_share2_reg ;
assign x1x3x4x7_second_share =      x1_share2_reg & x3x4x7_second_share ^    x3_share2_reg & x1x4x7_second_share ^    x1x3_share2_reg  & x4x7_second_share ^     x4_share2_reg  & x1x3x7_subscript0_share2_reg ^ x7_share2_reg  & x1x3x4_subscript0_share2_reg ^    x4x7_share2_reg  & x1x3_subscript0_share2_reg ^x1x3x4x7_subscript0_share2_reg ;
assign x1x3x5x6_second_share =      x1_share2_reg & x3x5x6_second_share ^    x3_share2_reg & x1x5x6_second_share ^    x1x3_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x1x3x6_subscript0_share2_reg ^ x6_share2_reg  & x1x3x5_subscript0_share2_reg ^    x5x6_share2_reg  & x1x3_subscript0_share2_reg ^x1x3x5x6_subscript0_share2_reg ;
assign x1x3x5x7_second_share =      x1_share2_reg & x3x5x7_second_share ^    x3_share2_reg & x1x5x7_second_share ^    x1x3_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x1x3x7_subscript0_share2_reg ^ x7_share2_reg  & x1x3x5_subscript0_share2_reg ^    x5x7_share2_reg  & x1x3_subscript0_share2_reg ^x1x3x5x7_subscript0_share2_reg ;
assign x1x3x6x7_second_share =      x1_share2_reg & x3x6x7_second_share ^    x3_share2_reg & x1x6x7_second_share ^    x1x3_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x1x3x7_subscript0_share2_reg ^ x7_share2_reg  & x1x3x6_subscript0_share2_reg ^    x6x7_share2_reg  & x1x3_subscript0_share2_reg ^x1x3x6x7_subscript0_share2_reg ;
assign x1x4x5x6_second_share =      x1_share2_reg & x4x5x6_second_share ^    x4_share2_reg & x1x5x6_second_share ^    x1x4_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x1x4x6_subscript0_share2_reg ^ x6_share2_reg  & x1x4x5_subscript0_share2_reg ^    x5x6_share2_reg  & x1x4_subscript0_share2_reg ^x1x4x5x6_subscript0_share2_reg ;
assign x1x4x5x7_second_share =      x1_share2_reg & x4x5x7_second_share ^    x4_share2_reg & x1x5x7_second_share ^    x1x4_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x1x4x7_subscript0_share2_reg ^ x7_share2_reg  & x1x4x5_subscript0_share2_reg ^    x5x7_share2_reg  & x1x4_subscript0_share2_reg ^x1x4x5x7_subscript0_share2_reg ;
assign x1x4x6x7_second_share =      x1_share2_reg & x4x6x7_second_share ^    x4_share2_reg & x1x6x7_second_share ^    x1x4_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x1x4x7_subscript0_share2_reg ^ x7_share2_reg  & x1x4x6_subscript0_share2_reg ^    x6x7_share2_reg  & x1x4_subscript0_share2_reg ^x1x4x6x7_subscript0_share2_reg ;
assign x1x5x6x7_second_share =      x1_share2_reg & x5x6x7_second_share ^    x5_share2_reg & x1x6x7_second_share ^    x1x5_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x1x5x7_subscript0_share2_reg ^ x7_share2_reg  & x1x5x6_subscript0_share2_reg ^    x6x7_share2_reg  & x1x5_subscript0_share2_reg ^x1x5x6x7_subscript0_share2_reg ;
assign x2x3x4x5_second_share =      x2_share2_reg & x3x4x5_second_share ^    x3_share2_reg & x2x4x5_second_share ^    x2x3_share2_reg  & x4x5_second_share ^     x4_share2_reg  & x2x3x5_subscript0_share2_reg ^ x5_share2_reg  & x2x3x4_subscript0_share2_reg ^    x4x5_share2_reg  & x2x3_subscript0_share2_reg ^x2x3x4x5_subscript0_share2_reg ;
assign x2x3x4x6_second_share =      x2_share2_reg & x3x4x6_second_share ^    x3_share2_reg & x2x4x6_second_share ^    x2x3_share2_reg  & x4x6_second_share ^     x4_share2_reg  & x2x3x6_subscript0_share2_reg ^ x6_share2_reg  & x2x3x4_subscript0_share2_reg ^    x4x6_share2_reg  & x2x3_subscript0_share2_reg ^x2x3x4x6_subscript0_share2_reg ;
assign x2x3x4x7_second_share =      x2_share2_reg & x3x4x7_second_share ^    x3_share2_reg & x2x4x7_second_share ^    x2x3_share2_reg  & x4x7_second_share ^     x4_share2_reg  & x2x3x7_subscript0_share2_reg ^ x7_share2_reg  & x2x3x4_subscript0_share2_reg ^    x4x7_share2_reg  & x2x3_subscript0_share2_reg ^x2x3x4x7_subscript0_share2_reg ;
assign x2x3x5x6_second_share =      x2_share2_reg & x3x5x6_second_share ^    x3_share2_reg & x2x5x6_second_share ^    x2x3_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x2x3x6_subscript0_share2_reg ^ x6_share2_reg  & x2x3x5_subscript0_share2_reg ^    x5x6_share2_reg  & x2x3_subscript0_share2_reg ^x2x3x5x6_subscript0_share2_reg ;
assign x2x3x5x7_second_share =      x2_share2_reg & x3x5x7_second_share ^    x3_share2_reg & x2x5x7_second_share ^    x2x3_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x2x3x7_subscript0_share2_reg ^ x7_share2_reg  & x2x3x5_subscript0_share2_reg ^    x5x7_share2_reg  & x2x3_subscript0_share2_reg ^x2x3x5x7_subscript0_share2_reg ;
assign x2x3x6x7_second_share =      x2_share2_reg & x3x6x7_second_share ^    x3_share2_reg & x2x6x7_second_share ^    x2x3_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x2x3x7_subscript0_share2_reg ^ x7_share2_reg  & x2x3x6_subscript0_share2_reg ^    x6x7_share2_reg  & x2x3_subscript0_share2_reg ^x2x3x6x7_subscript0_share2_reg ;
assign x2x4x5x6_second_share =      x2_share2_reg & x4x5x6_second_share ^    x4_share2_reg & x2x5x6_second_share ^    x2x4_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x2x4x6_subscript0_share2_reg ^ x6_share2_reg  & x2x4x5_subscript0_share2_reg ^    x5x6_share2_reg  & x2x4_subscript0_share2_reg ^x2x4x5x6_subscript0_share2_reg ;
assign x2x4x5x7_second_share =      x2_share2_reg & x4x5x7_second_share ^    x4_share2_reg & x2x5x7_second_share ^    x2x4_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x2x4x7_subscript0_share2_reg ^ x7_share2_reg  & x2x4x5_subscript0_share2_reg ^    x5x7_share2_reg  & x2x4_subscript0_share2_reg ^x2x4x5x7_subscript0_share2_reg ;
assign x2x4x6x7_second_share =      x2_share2_reg & x4x6x7_second_share ^    x4_share2_reg & x2x6x7_second_share ^    x2x4_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x2x4x7_subscript0_share2_reg ^ x7_share2_reg  & x2x4x6_subscript0_share2_reg ^    x6x7_share2_reg  & x2x4_subscript0_share2_reg ^x2x4x6x7_subscript0_share2_reg ;
assign x2x5x6x7_second_share =      x2_share2_reg & x5x6x7_second_share ^    x5_share2_reg & x2x6x7_second_share ^    x2x5_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x2x5x7_subscript0_share2_reg ^ x7_share2_reg  & x2x5x6_subscript0_share2_reg ^    x6x7_share2_reg  & x2x5_subscript0_share2_reg ^x2x5x6x7_subscript0_share2_reg ;
assign x3x4x5x6_second_share =      x3_share2_reg & x4x5x6_second_share ^    x4_share2_reg & x3x5x6_second_share ^    x3x4_share2_reg  & x5x6_second_share ^     x5_share2_reg  & x3x4x6_subscript0_share2_reg ^ x6_share2_reg  & x3x4x5_subscript0_share2_reg ^    x5x6_share2_reg  & x3x4_subscript0_share2_reg ^x3x4x5x6_subscript0_share2_reg ;
assign x3x4x5x7_second_share =      x3_share2_reg & x4x5x7_second_share ^    x4_share2_reg & x3x5x7_second_share ^    x3x4_share2_reg  & x5x7_second_share ^     x5_share2_reg  & x3x4x7_subscript0_share2_reg ^ x7_share2_reg  & x3x4x5_subscript0_share2_reg ^    x5x7_share2_reg  & x3x4_subscript0_share2_reg ^x3x4x5x7_subscript0_share2_reg ;
assign x3x4x6x7_second_share =      x3_share2_reg & x4x6x7_second_share ^    x4_share2_reg & x3x6x7_second_share ^    x3x4_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x3x4x7_subscript0_share2_reg ^ x7_share2_reg  & x3x4x6_subscript0_share2_reg ^    x6x7_share2_reg  & x3x4_subscript0_share2_reg ^x3x4x6x7_subscript0_share2_reg ;
assign x3x5x6x7_second_share =      x3_share2_reg & x5x6x7_second_share ^    x5_share2_reg & x3x6x7_second_share ^    x3x5_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x3x5x7_subscript0_share2_reg ^ x7_share2_reg  & x3x5x6_subscript0_share2_reg ^    x6x7_share2_reg  & x3x5_subscript0_share2_reg ^x3x5x6x7_subscript0_share2_reg ;
assign x4x5x6x7_second_share =      x4_share2_reg & x5x6x7_second_share ^    x5_share2_reg & x4x6x7_second_share ^    x4x5_share2_reg  & x6x7_second_share ^     x6_share2_reg  & x4x5x7_subscript0_share2_reg ^ x7_share2_reg  & x4x5x6_subscript0_share2_reg ^    x6x7_share2_reg  & x4x5_subscript0_share2_reg ^x4x5x6x7_subscript0_share2_reg ;


// second share of Degree-5 terms

assign x0x1x2x3x4_second_share =x0_share2_reg & x1x2x3x4_second_share ^ x1_share2_reg & x0x2x3x4_second_share ^ x0x1_share2_reg & x2x3x4_second_share ^ x2x3x4_share2_reg & x0x1_subscript0_share2_reg ^x2x3_share2_reg & x0x1x4_subscript0_share2_reg ^x2x4_share2_reg & x0x1x3_subscript0_share2_reg ^x3x4_share2_reg & x0x1x2_subscript0_share2_reg ^x4_share2_reg & x0x1x2x3_subscript0_share2_reg ^x3_share2_reg & x0x1x2x4_subscript0_share2_reg ^x2_share2_reg & x0x1x3x4_subscript0_share2_reg ^x0x1x2x3x4_subscript0_share2_reg ;
assign x0x1x2x3x5_second_share =x0_share2_reg & x1x2x3x5_second_share ^ x1_share2_reg & x0x2x3x5_second_share ^ x0x1_share2_reg & x2x3x5_second_share ^ x2x3x5_share2_reg & x0x1_subscript0_share2_reg ^x2x3_share2_reg & x0x1x5_subscript0_share2_reg ^x2x5_share2_reg & x0x1x3_subscript0_share2_reg ^x3x5_share2_reg & x0x1x2_subscript0_share2_reg ^x5_share2_reg & x0x1x2x3_subscript0_share2_reg ^x3_share2_reg & x0x1x2x5_subscript0_share2_reg ^x2_share2_reg & x0x1x3x5_subscript0_share2_reg ^x0x1x2x3x5_subscript0_share2_reg ;
assign x0x1x2x3x6_second_share =x0_share2_reg & x1x2x3x6_second_share ^ x1_share2_reg & x0x2x3x6_second_share ^ x0x1_share2_reg & x2x3x6_second_share ^ x2x3x6_share2_reg & x0x1_subscript0_share2_reg ^x2x3_share2_reg & x0x1x6_subscript0_share2_reg ^x2x6_share2_reg & x0x1x3_subscript0_share2_reg ^x3x6_share2_reg & x0x1x2_subscript0_share2_reg ^x6_share2_reg & x0x1x2x3_subscript0_share2_reg ^x3_share2_reg & x0x1x2x6_subscript0_share2_reg ^x2_share2_reg & x0x1x3x6_subscript0_share2_reg ^x0x1x2x3x6_subscript0_share2_reg ;
assign x0x1x2x3x7_second_share =x0_share2_reg & x1x2x3x7_second_share ^ x1_share2_reg & x0x2x3x7_second_share ^ x0x1_share2_reg & x2x3x7_second_share ^ x2x3x7_share2_reg & x0x1_subscript0_share2_reg ^x2x3_share2_reg & x0x1x7_subscript0_share2_reg ^x2x7_share2_reg & x0x1x3_subscript0_share2_reg ^x3x7_share2_reg & x0x1x2_subscript0_share2_reg ^x7_share2_reg & x0x1x2x3_subscript0_share2_reg ^x3_share2_reg & x0x1x2x7_subscript0_share2_reg ^x2_share2_reg & x0x1x3x7_subscript0_share2_reg ^x0x1x2x3x7_subscript0_share2_reg ;
assign x0x1x2x4x5_second_share =x0_share2_reg & x1x2x4x5_second_share ^ x1_share2_reg & x0x2x4x5_second_share ^ x0x1_share2_reg & x2x4x5_second_share ^ x2x4x5_share2_reg & x0x1_subscript0_share2_reg ^x2x4_share2_reg & x0x1x5_subscript0_share2_reg ^x2x5_share2_reg & x0x1x4_subscript0_share2_reg ^x4x5_share2_reg & x0x1x2_subscript0_share2_reg ^x5_share2_reg & x0x1x2x4_subscript0_share2_reg ^x4_share2_reg & x0x1x2x5_subscript0_share2_reg ^x2_share2_reg & x0x1x4x5_subscript0_share2_reg ^x0x1x2x4x5_subscript0_share2_reg ;
assign x0x1x2x4x6_second_share =x0_share2_reg & x1x2x4x6_second_share ^ x1_share2_reg & x0x2x4x6_second_share ^ x0x1_share2_reg & x2x4x6_second_share ^ x2x4x6_share2_reg & x0x1_subscript0_share2_reg ^x2x4_share2_reg & x0x1x6_subscript0_share2_reg ^x2x6_share2_reg & x0x1x4_subscript0_share2_reg ^x4x6_share2_reg & x0x1x2_subscript0_share2_reg ^x6_share2_reg & x0x1x2x4_subscript0_share2_reg ^x4_share2_reg & x0x1x2x6_subscript0_share2_reg ^x2_share2_reg & x0x1x4x6_subscript0_share2_reg ^x0x1x2x4x6_subscript0_share2_reg ;
assign x0x1x2x4x7_second_share =x0_share2_reg & x1x2x4x7_second_share ^ x1_share2_reg & x0x2x4x7_second_share ^ x0x1_share2_reg & x2x4x7_second_share ^ x2x4x7_share2_reg & x0x1_subscript0_share2_reg ^x2x4_share2_reg & x0x1x7_subscript0_share2_reg ^x2x7_share2_reg & x0x1x4_subscript0_share2_reg ^x4x7_share2_reg & x0x1x2_subscript0_share2_reg ^x7_share2_reg & x0x1x2x4_subscript0_share2_reg ^x4_share2_reg & x0x1x2x7_subscript0_share2_reg ^x2_share2_reg & x0x1x4x7_subscript0_share2_reg ^x0x1x2x4x7_subscript0_share2_reg ;
assign x0x1x2x5x6_second_share =x0_share2_reg & x1x2x5x6_second_share ^ x1_share2_reg & x0x2x5x6_second_share ^ x0x1_share2_reg & x2x5x6_second_share ^ x2x5x6_share2_reg & x0x1_subscript0_share2_reg ^x2x5_share2_reg & x0x1x6_subscript0_share2_reg ^x2x6_share2_reg & x0x1x5_subscript0_share2_reg ^x5x6_share2_reg & x0x1x2_subscript0_share2_reg ^x6_share2_reg & x0x1x2x5_subscript0_share2_reg ^x5_share2_reg & x0x1x2x6_subscript0_share2_reg ^x2_share2_reg & x0x1x5x6_subscript0_share2_reg ^x0x1x2x5x6_subscript0_share2_reg ;
assign x0x1x2x5x7_second_share =x0_share2_reg & x1x2x5x7_second_share ^ x1_share2_reg & x0x2x5x7_second_share ^ x0x1_share2_reg & x2x5x7_second_share ^ x2x5x7_share2_reg & x0x1_subscript0_share2_reg ^x2x5_share2_reg & x0x1x7_subscript0_share2_reg ^x2x7_share2_reg & x0x1x5_subscript0_share2_reg ^x5x7_share2_reg & x0x1x2_subscript0_share2_reg ^x7_share2_reg & x0x1x2x5_subscript0_share2_reg ^x5_share2_reg & x0x1x2x7_subscript0_share2_reg ^x2_share2_reg & x0x1x5x7_subscript0_share2_reg ^x0x1x2x5x7_subscript0_share2_reg ;
assign x0x1x2x6x7_second_share =x0_share2_reg & x1x2x6x7_second_share ^ x1_share2_reg & x0x2x6x7_second_share ^ x0x1_share2_reg & x2x6x7_second_share ^ x2x6x7_share2_reg & x0x1_subscript0_share2_reg ^x2x6_share2_reg & x0x1x7_subscript0_share2_reg ^x2x7_share2_reg & x0x1x6_subscript0_share2_reg ^x6x7_share2_reg & x0x1x2_subscript0_share2_reg ^x7_share2_reg & x0x1x2x6_subscript0_share2_reg ^x6_share2_reg & x0x1x2x7_subscript0_share2_reg ^x2_share2_reg & x0x1x6x7_subscript0_share2_reg ^x0x1x2x6x7_subscript0_share2_reg ;
assign x0x1x3x4x5_second_share =x0_share2_reg & x1x3x4x5_second_share ^ x1_share2_reg & x0x3x4x5_second_share ^ x0x1_share2_reg & x3x4x5_second_share ^ x3x4x5_share2_reg & x0x1_subscript0_share2_reg ^x3x4_share2_reg & x0x1x5_subscript0_share2_reg ^x3x5_share2_reg & x0x1x4_subscript0_share2_reg ^x4x5_share2_reg & x0x1x3_subscript0_share2_reg ^x5_share2_reg & x0x1x3x4_subscript0_share2_reg ^x4_share2_reg & x0x1x3x5_subscript0_share2_reg ^x3_share2_reg & x0x1x4x5_subscript0_share2_reg ^x0x1x3x4x5_subscript0_share2_reg ;
assign x0x1x3x4x6_second_share =x0_share2_reg & x1x3x4x6_second_share ^ x1_share2_reg & x0x3x4x6_second_share ^ x0x1_share2_reg & x3x4x6_second_share ^ x3x4x6_share2_reg & x0x1_subscript0_share2_reg ^x3x4_share2_reg & x0x1x6_subscript0_share2_reg ^x3x6_share2_reg & x0x1x4_subscript0_share2_reg ^x4x6_share2_reg & x0x1x3_subscript0_share2_reg ^x6_share2_reg & x0x1x3x4_subscript0_share2_reg ^x4_share2_reg & x0x1x3x6_subscript0_share2_reg ^x3_share2_reg & x0x1x4x6_subscript0_share2_reg ^x0x1x3x4x6_subscript0_share2_reg ;
assign x0x1x3x4x7_second_share =x0_share2_reg & x1x3x4x7_second_share ^ x1_share2_reg & x0x3x4x7_second_share ^ x0x1_share2_reg & x3x4x7_second_share ^ x3x4x7_share2_reg & x0x1_subscript0_share2_reg ^x3x4_share2_reg & x0x1x7_subscript0_share2_reg ^x3x7_share2_reg & x0x1x4_subscript0_share2_reg ^x4x7_share2_reg & x0x1x3_subscript0_share2_reg ^x7_share2_reg & x0x1x3x4_subscript0_share2_reg ^x4_share2_reg & x0x1x3x7_subscript0_share2_reg ^x3_share2_reg & x0x1x4x7_subscript0_share2_reg ^x0x1x3x4x7_subscript0_share2_reg ;
assign x0x1x3x5x6_second_share =x0_share2_reg & x1x3x5x6_second_share ^ x1_share2_reg & x0x3x5x6_second_share ^ x0x1_share2_reg & x3x5x6_second_share ^ x3x5x6_share2_reg & x0x1_subscript0_share2_reg ^x3x5_share2_reg & x0x1x6_subscript0_share2_reg ^x3x6_share2_reg & x0x1x5_subscript0_share2_reg ^x5x6_share2_reg & x0x1x3_subscript0_share2_reg ^x6_share2_reg & x0x1x3x5_subscript0_share2_reg ^x5_share2_reg & x0x1x3x6_subscript0_share2_reg ^x3_share2_reg & x0x1x5x6_subscript0_share2_reg ^x0x1x3x5x6_subscript0_share2_reg ;
assign x0x1x3x5x7_second_share =x0_share2_reg & x1x3x5x7_second_share ^ x1_share2_reg & x0x3x5x7_second_share ^ x0x1_share2_reg & x3x5x7_second_share ^ x3x5x7_share2_reg & x0x1_subscript0_share2_reg ^x3x5_share2_reg & x0x1x7_subscript0_share2_reg ^x3x7_share2_reg & x0x1x5_subscript0_share2_reg ^x5x7_share2_reg & x0x1x3_subscript0_share2_reg ^x7_share2_reg & x0x1x3x5_subscript0_share2_reg ^x5_share2_reg & x0x1x3x7_subscript0_share2_reg ^x3_share2_reg & x0x1x5x7_subscript0_share2_reg ^x0x1x3x5x7_subscript0_share2_reg ;
assign x0x1x3x6x7_second_share =x0_share2_reg & x1x3x6x7_second_share ^ x1_share2_reg & x0x3x6x7_second_share ^ x0x1_share2_reg & x3x6x7_second_share ^ x3x6x7_share2_reg & x0x1_subscript0_share2_reg ^x3x6_share2_reg & x0x1x7_subscript0_share2_reg ^x3x7_share2_reg & x0x1x6_subscript0_share2_reg ^x6x7_share2_reg & x0x1x3_subscript0_share2_reg ^x7_share2_reg & x0x1x3x6_subscript0_share2_reg ^x6_share2_reg & x0x1x3x7_subscript0_share2_reg ^x3_share2_reg & x0x1x6x7_subscript0_share2_reg ^x0x1x3x6x7_subscript0_share2_reg ;
assign x0x1x4x5x6_second_share =x0_share2_reg & x1x4x5x6_second_share ^ x1_share2_reg & x0x4x5x6_second_share ^ x0x1_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x0x1_subscript0_share2_reg ^x4x5_share2_reg & x0x1x6_subscript0_share2_reg ^x4x6_share2_reg & x0x1x5_subscript0_share2_reg ^x5x6_share2_reg & x0x1x4_subscript0_share2_reg ^x6_share2_reg & x0x1x4x5_subscript0_share2_reg ^x5_share2_reg & x0x1x4x6_subscript0_share2_reg ^x4_share2_reg & x0x1x5x6_subscript0_share2_reg ^x0x1x4x5x6_subscript0_share2_reg ;
assign x0x1x4x5x7_second_share =x0_share2_reg & x1x4x5x7_second_share ^ x1_share2_reg & x0x4x5x7_second_share ^ x0x1_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x0x1_subscript0_share2_reg ^x4x5_share2_reg & x0x1x7_subscript0_share2_reg ^x4x7_share2_reg & x0x1x5_subscript0_share2_reg ^x5x7_share2_reg & x0x1x4_subscript0_share2_reg ^x7_share2_reg & x0x1x4x5_subscript0_share2_reg ^x5_share2_reg & x0x1x4x7_subscript0_share2_reg ^x4_share2_reg & x0x1x5x7_subscript0_share2_reg ^x0x1x4x5x7_subscript0_share2_reg ;
assign x0x1x4x6x7_second_share =x0_share2_reg & x1x4x6x7_second_share ^ x1_share2_reg & x0x4x6x7_second_share ^ x0x1_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x0x1_subscript0_share2_reg ^x4x6_share2_reg & x0x1x7_subscript0_share2_reg ^x4x7_share2_reg & x0x1x6_subscript0_share2_reg ^x6x7_share2_reg & x0x1x4_subscript0_share2_reg ^x7_share2_reg & x0x1x4x6_subscript0_share2_reg ^x6_share2_reg & x0x1x4x7_subscript0_share2_reg ^x4_share2_reg & x0x1x6x7_subscript0_share2_reg ^x0x1x4x6x7_subscript0_share2_reg ;
assign x0x1x5x6x7_second_share =x0_share2_reg & x1x5x6x7_second_share ^ x1_share2_reg & x0x5x6x7_second_share ^ x0x1_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x1_subscript0_share2_reg ^x5x6_share2_reg & x0x1x7_subscript0_share2_reg ^x5x7_share2_reg & x0x1x6_subscript0_share2_reg ^x6x7_share2_reg & x0x1x5_subscript0_share2_reg ^x7_share2_reg & x0x1x5x6_subscript0_share2_reg ^x6_share2_reg & x0x1x5x7_subscript0_share2_reg ^x5_share2_reg & x0x1x6x7_subscript0_share2_reg ^x0x1x5x6x7_subscript0_share2_reg ;
assign x0x2x3x4x5_second_share =x0_share2_reg & x2x3x4x5_second_share ^ x2_share2_reg & x0x3x4x5_second_share ^ x0x2_share2_reg & x3x4x5_second_share ^ x3x4x5_share2_reg & x0x2_subscript0_share2_reg ^x3x4_share2_reg & x0x2x5_subscript0_share2_reg ^x3x5_share2_reg & x0x2x4_subscript0_share2_reg ^x4x5_share2_reg & x0x2x3_subscript0_share2_reg ^x5_share2_reg & x0x2x3x4_subscript0_share2_reg ^x4_share2_reg & x0x2x3x5_subscript0_share2_reg ^x3_share2_reg & x0x2x4x5_subscript0_share2_reg ^x0x2x3x4x5_subscript0_share2_reg ;
assign x0x2x3x4x6_second_share =x0_share2_reg & x2x3x4x6_second_share ^ x2_share2_reg & x0x3x4x6_second_share ^ x0x2_share2_reg & x3x4x6_second_share ^ x3x4x6_share2_reg & x0x2_subscript0_share2_reg ^x3x4_share2_reg & x0x2x6_subscript0_share2_reg ^x3x6_share2_reg & x0x2x4_subscript0_share2_reg ^x4x6_share2_reg & x0x2x3_subscript0_share2_reg ^x6_share2_reg & x0x2x3x4_subscript0_share2_reg ^x4_share2_reg & x0x2x3x6_subscript0_share2_reg ^x3_share2_reg & x0x2x4x6_subscript0_share2_reg ^x0x2x3x4x6_subscript0_share2_reg ;
assign x0x2x3x4x7_second_share =x0_share2_reg & x2x3x4x7_second_share ^ x2_share2_reg & x0x3x4x7_second_share ^ x0x2_share2_reg & x3x4x7_second_share ^ x3x4x7_share2_reg & x0x2_subscript0_share2_reg ^x3x4_share2_reg & x0x2x7_subscript0_share2_reg ^x3x7_share2_reg & x0x2x4_subscript0_share2_reg ^x4x7_share2_reg & x0x2x3_subscript0_share2_reg ^x7_share2_reg & x0x2x3x4_subscript0_share2_reg ^x4_share2_reg & x0x2x3x7_subscript0_share2_reg ^x3_share2_reg & x0x2x4x7_subscript0_share2_reg ^x0x2x3x4x7_subscript0_share2_reg ;
assign x0x2x3x5x6_second_share =x0_share2_reg & x2x3x5x6_second_share ^ x2_share2_reg & x0x3x5x6_second_share ^ x0x2_share2_reg & x3x5x6_second_share ^ x3x5x6_share2_reg & x0x2_subscript0_share2_reg ^x3x5_share2_reg & x0x2x6_subscript0_share2_reg ^x3x6_share2_reg & x0x2x5_subscript0_share2_reg ^x5x6_share2_reg & x0x2x3_subscript0_share2_reg ^x6_share2_reg & x0x2x3x5_subscript0_share2_reg ^x5_share2_reg & x0x2x3x6_subscript0_share2_reg ^x3_share2_reg & x0x2x5x6_subscript0_share2_reg ^x0x2x3x5x6_subscript0_share2_reg ;
assign x0x2x3x5x7_second_share =x0_share2_reg & x2x3x5x7_second_share ^ x2_share2_reg & x0x3x5x7_second_share ^ x0x2_share2_reg & x3x5x7_second_share ^ x3x5x7_share2_reg & x0x2_subscript0_share2_reg ^x3x5_share2_reg & x0x2x7_subscript0_share2_reg ^x3x7_share2_reg & x0x2x5_subscript0_share2_reg ^x5x7_share2_reg & x0x2x3_subscript0_share2_reg ^x7_share2_reg & x0x2x3x5_subscript0_share2_reg ^x5_share2_reg & x0x2x3x7_subscript0_share2_reg ^x3_share2_reg & x0x2x5x7_subscript0_share2_reg ^x0x2x3x5x7_subscript0_share2_reg ;
assign x0x2x3x6x7_second_share =x0_share2_reg & x2x3x6x7_second_share ^ x2_share2_reg & x0x3x6x7_second_share ^ x0x2_share2_reg & x3x6x7_second_share ^ x3x6x7_share2_reg & x0x2_subscript0_share2_reg ^x3x6_share2_reg & x0x2x7_subscript0_share2_reg ^x3x7_share2_reg & x0x2x6_subscript0_share2_reg ^x6x7_share2_reg & x0x2x3_subscript0_share2_reg ^x7_share2_reg & x0x2x3x6_subscript0_share2_reg ^x6_share2_reg & x0x2x3x7_subscript0_share2_reg ^x3_share2_reg & x0x2x6x7_subscript0_share2_reg ^x0x2x3x6x7_subscript0_share2_reg ;
assign x0x2x4x5x6_second_share =x0_share2_reg & x2x4x5x6_second_share ^ x2_share2_reg & x0x4x5x6_second_share ^ x0x2_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x0x2_subscript0_share2_reg ^x4x5_share2_reg & x0x2x6_subscript0_share2_reg ^x4x6_share2_reg & x0x2x5_subscript0_share2_reg ^x5x6_share2_reg & x0x2x4_subscript0_share2_reg ^x6_share2_reg & x0x2x4x5_subscript0_share2_reg ^x5_share2_reg & x0x2x4x6_subscript0_share2_reg ^x4_share2_reg & x0x2x5x6_subscript0_share2_reg ^x0x2x4x5x6_subscript0_share2_reg ;
assign x0x2x4x5x7_second_share =x0_share2_reg & x2x4x5x7_second_share ^ x2_share2_reg & x0x4x5x7_second_share ^ x0x2_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x0x2_subscript0_share2_reg ^x4x5_share2_reg & x0x2x7_subscript0_share2_reg ^x4x7_share2_reg & x0x2x5_subscript0_share2_reg ^x5x7_share2_reg & x0x2x4_subscript0_share2_reg ^x7_share2_reg & x0x2x4x5_subscript0_share2_reg ^x5_share2_reg & x0x2x4x7_subscript0_share2_reg ^x4_share2_reg & x0x2x5x7_subscript0_share2_reg ^x0x2x4x5x7_subscript0_share2_reg ;
assign x0x2x4x6x7_second_share =x0_share2_reg & x2x4x6x7_second_share ^ x2_share2_reg & x0x4x6x7_second_share ^ x0x2_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x0x2_subscript0_share2_reg ^x4x6_share2_reg & x0x2x7_subscript0_share2_reg ^x4x7_share2_reg & x0x2x6_subscript0_share2_reg ^x6x7_share2_reg & x0x2x4_subscript0_share2_reg ^x7_share2_reg & x0x2x4x6_subscript0_share2_reg ^x6_share2_reg & x0x2x4x7_subscript0_share2_reg ^x4_share2_reg & x0x2x6x7_subscript0_share2_reg ^x0x2x4x6x7_subscript0_share2_reg ;
assign x0x2x5x6x7_second_share =x0_share2_reg & x2x5x6x7_second_share ^ x2_share2_reg & x0x5x6x7_second_share ^ x0x2_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x2_subscript0_share2_reg ^x5x6_share2_reg & x0x2x7_subscript0_share2_reg ^x5x7_share2_reg & x0x2x6_subscript0_share2_reg ^x6x7_share2_reg & x0x2x5_subscript0_share2_reg ^x7_share2_reg & x0x2x5x6_subscript0_share2_reg ^x6_share2_reg & x0x2x5x7_subscript0_share2_reg ^x5_share2_reg & x0x2x6x7_subscript0_share2_reg ^x0x2x5x6x7_subscript0_share2_reg ;
assign x0x3x4x5x6_second_share =x0_share2_reg & x3x4x5x6_second_share ^ x3_share2_reg & x0x4x5x6_second_share ^ x0x3_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x0x3_subscript0_share2_reg ^x4x5_share2_reg & x0x3x6_subscript0_share2_reg ^x4x6_share2_reg & x0x3x5_subscript0_share2_reg ^x5x6_share2_reg & x0x3x4_subscript0_share2_reg ^x6_share2_reg & x0x3x4x5_subscript0_share2_reg ^x5_share2_reg & x0x3x4x6_subscript0_share2_reg ^x4_share2_reg & x0x3x5x6_subscript0_share2_reg ^x0x3x4x5x6_subscript0_share2_reg ;
assign x0x3x4x5x7_second_share =x0_share2_reg & x3x4x5x7_second_share ^ x3_share2_reg & x0x4x5x7_second_share ^ x0x3_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x0x3_subscript0_share2_reg ^x4x5_share2_reg & x0x3x7_subscript0_share2_reg ^x4x7_share2_reg & x0x3x5_subscript0_share2_reg ^x5x7_share2_reg & x0x3x4_subscript0_share2_reg ^x7_share2_reg & x0x3x4x5_subscript0_share2_reg ^x5_share2_reg & x0x3x4x7_subscript0_share2_reg ^x4_share2_reg & x0x3x5x7_subscript0_share2_reg ^x0x3x4x5x7_subscript0_share2_reg ;
assign x0x3x4x6x7_second_share =x0_share2_reg & x3x4x6x7_second_share ^ x3_share2_reg & x0x4x6x7_second_share ^ x0x3_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x0x3_subscript0_share2_reg ^x4x6_share2_reg & x0x3x7_subscript0_share2_reg ^x4x7_share2_reg & x0x3x6_subscript0_share2_reg ^x6x7_share2_reg & x0x3x4_subscript0_share2_reg ^x7_share2_reg & x0x3x4x6_subscript0_share2_reg ^x6_share2_reg & x0x3x4x7_subscript0_share2_reg ^x4_share2_reg & x0x3x6x7_subscript0_share2_reg ^x0x3x4x6x7_subscript0_share2_reg ;
assign x0x3x5x6x7_second_share =x0_share2_reg & x3x5x6x7_second_share ^ x3_share2_reg & x0x5x6x7_second_share ^ x0x3_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x3_subscript0_share2_reg ^x5x6_share2_reg & x0x3x7_subscript0_share2_reg ^x5x7_share2_reg & x0x3x6_subscript0_share2_reg ^x6x7_share2_reg & x0x3x5_subscript0_share2_reg ^x7_share2_reg & x0x3x5x6_subscript0_share2_reg ^x6_share2_reg & x0x3x5x7_subscript0_share2_reg ^x5_share2_reg & x0x3x6x7_subscript0_share2_reg ^x0x3x5x6x7_subscript0_share2_reg ;
assign x0x4x5x6x7_second_share =x0_share2_reg & x4x5x6x7_second_share ^ x4_share2_reg & x0x5x6x7_second_share ^ x0x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x4_subscript0_share2_reg ^x5x6_share2_reg & x0x4x7_subscript0_share2_reg ^x5x7_share2_reg & x0x4x6_subscript0_share2_reg ^x6x7_share2_reg & x0x4x5_subscript0_share2_reg ^x7_share2_reg & x0x4x5x6_subscript0_share2_reg ^x6_share2_reg & x0x4x5x7_subscript0_share2_reg ^x5_share2_reg & x0x4x6x7_subscript0_share2_reg ^x0x4x5x6x7_subscript0_share2_reg ;
assign x1x2x3x4x5_second_share =x1_share2_reg & x2x3x4x5_second_share ^ x2_share2_reg & x1x3x4x5_second_share ^ x1x2_share2_reg & x3x4x5_second_share ^ x3x4x5_share2_reg & x1x2_subscript0_share2_reg ^x3x4_share2_reg & x1x2x5_subscript0_share2_reg ^x3x5_share2_reg & x1x2x4_subscript0_share2_reg ^x4x5_share2_reg & x1x2x3_subscript0_share2_reg ^x5_share2_reg & x1x2x3x4_subscript0_share2_reg ^x4_share2_reg & x1x2x3x5_subscript0_share2_reg ^x3_share2_reg & x1x2x4x5_subscript0_share2_reg ^x1x2x3x4x5_subscript0_share2_reg ;
assign x1x2x3x4x6_second_share =x1_share2_reg & x2x3x4x6_second_share ^ x2_share2_reg & x1x3x4x6_second_share ^ x1x2_share2_reg & x3x4x6_second_share ^ x3x4x6_share2_reg & x1x2_subscript0_share2_reg ^x3x4_share2_reg & x1x2x6_subscript0_share2_reg ^x3x6_share2_reg & x1x2x4_subscript0_share2_reg ^x4x6_share2_reg & x1x2x3_subscript0_share2_reg ^x6_share2_reg & x1x2x3x4_subscript0_share2_reg ^x4_share2_reg & x1x2x3x6_subscript0_share2_reg ^x3_share2_reg & x1x2x4x6_subscript0_share2_reg ^x1x2x3x4x6_subscript0_share2_reg ;
assign x1x2x3x4x7_second_share =x1_share2_reg & x2x3x4x7_second_share ^ x2_share2_reg & x1x3x4x7_second_share ^ x1x2_share2_reg & x3x4x7_second_share ^ x3x4x7_share2_reg & x1x2_subscript0_share2_reg ^x3x4_share2_reg & x1x2x7_subscript0_share2_reg ^x3x7_share2_reg & x1x2x4_subscript0_share2_reg ^x4x7_share2_reg & x1x2x3_subscript0_share2_reg ^x7_share2_reg & x1x2x3x4_subscript0_share2_reg ^x4_share2_reg & x1x2x3x7_subscript0_share2_reg ^x3_share2_reg & x1x2x4x7_subscript0_share2_reg ^x1x2x3x4x7_subscript0_share2_reg ;
assign x1x2x3x5x6_second_share =x1_share2_reg & x2x3x5x6_second_share ^ x2_share2_reg & x1x3x5x6_second_share ^ x1x2_share2_reg & x3x5x6_second_share ^ x3x5x6_share2_reg & x1x2_subscript0_share2_reg ^x3x5_share2_reg & x1x2x6_subscript0_share2_reg ^x3x6_share2_reg & x1x2x5_subscript0_share2_reg ^x5x6_share2_reg & x1x2x3_subscript0_share2_reg ^x6_share2_reg & x1x2x3x5_subscript0_share2_reg ^x5_share2_reg & x1x2x3x6_subscript0_share2_reg ^x3_share2_reg & x1x2x5x6_subscript0_share2_reg ^x1x2x3x5x6_subscript0_share2_reg ;
assign x1x2x3x5x7_second_share =x1_share2_reg & x2x3x5x7_second_share ^ x2_share2_reg & x1x3x5x7_second_share ^ x1x2_share2_reg & x3x5x7_second_share ^ x3x5x7_share2_reg & x1x2_subscript0_share2_reg ^x3x5_share2_reg & x1x2x7_subscript0_share2_reg ^x3x7_share2_reg & x1x2x5_subscript0_share2_reg ^x5x7_share2_reg & x1x2x3_subscript0_share2_reg ^x7_share2_reg & x1x2x3x5_subscript0_share2_reg ^x5_share2_reg & x1x2x3x7_subscript0_share2_reg ^x3_share2_reg & x1x2x5x7_subscript0_share2_reg ^x1x2x3x5x7_subscript0_share2_reg ;
assign x1x2x3x6x7_second_share =x1_share2_reg & x2x3x6x7_second_share ^ x2_share2_reg & x1x3x6x7_second_share ^ x1x2_share2_reg & x3x6x7_second_share ^ x3x6x7_share2_reg & x1x2_subscript0_share2_reg ^x3x6_share2_reg & x1x2x7_subscript0_share2_reg ^x3x7_share2_reg & x1x2x6_subscript0_share2_reg ^x6x7_share2_reg & x1x2x3_subscript0_share2_reg ^x7_share2_reg & x1x2x3x6_subscript0_share2_reg ^x6_share2_reg & x1x2x3x7_subscript0_share2_reg ^x3_share2_reg & x1x2x6x7_subscript0_share2_reg ^x1x2x3x6x7_subscript0_share2_reg ;
assign x1x2x4x5x6_second_share =x1_share2_reg & x2x4x5x6_second_share ^ x2_share2_reg & x1x4x5x6_second_share ^ x1x2_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x1x2_subscript0_share2_reg ^x4x5_share2_reg & x1x2x6_subscript0_share2_reg ^x4x6_share2_reg & x1x2x5_subscript0_share2_reg ^x5x6_share2_reg & x1x2x4_subscript0_share2_reg ^x6_share2_reg & x1x2x4x5_subscript0_share2_reg ^x5_share2_reg & x1x2x4x6_subscript0_share2_reg ^x4_share2_reg & x1x2x5x6_subscript0_share2_reg ^x1x2x4x5x6_subscript0_share2_reg ;
assign x1x2x4x5x7_second_share =x1_share2_reg & x2x4x5x7_second_share ^ x2_share2_reg & x1x4x5x7_second_share ^ x1x2_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x1x2_subscript0_share2_reg ^x4x5_share2_reg & x1x2x7_subscript0_share2_reg ^x4x7_share2_reg & x1x2x5_subscript0_share2_reg ^x5x7_share2_reg & x1x2x4_subscript0_share2_reg ^x7_share2_reg & x1x2x4x5_subscript0_share2_reg ^x5_share2_reg & x1x2x4x7_subscript0_share2_reg ^x4_share2_reg & x1x2x5x7_subscript0_share2_reg ^x1x2x4x5x7_subscript0_share2_reg ;
assign x1x2x4x6x7_second_share =x1_share2_reg & x2x4x6x7_second_share ^ x2_share2_reg & x1x4x6x7_second_share ^ x1x2_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x1x2_subscript0_share2_reg ^x4x6_share2_reg & x1x2x7_subscript0_share2_reg ^x4x7_share2_reg & x1x2x6_subscript0_share2_reg ^x6x7_share2_reg & x1x2x4_subscript0_share2_reg ^x7_share2_reg & x1x2x4x6_subscript0_share2_reg ^x6_share2_reg & x1x2x4x7_subscript0_share2_reg ^x4_share2_reg & x1x2x6x7_subscript0_share2_reg ^x1x2x4x6x7_subscript0_share2_reg ;
assign x1x2x5x6x7_second_share =x1_share2_reg & x2x5x6x7_second_share ^ x2_share2_reg & x1x5x6x7_second_share ^ x1x2_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x1x2_subscript0_share2_reg ^x5x6_share2_reg & x1x2x7_subscript0_share2_reg ^x5x7_share2_reg & x1x2x6_subscript0_share2_reg ^x6x7_share2_reg & x1x2x5_subscript0_share2_reg ^x7_share2_reg & x1x2x5x6_subscript0_share2_reg ^x6_share2_reg & x1x2x5x7_subscript0_share2_reg ^x5_share2_reg & x1x2x6x7_subscript0_share2_reg ^x1x2x5x6x7_subscript0_share2_reg ;
assign x1x3x4x5x6_second_share =x1_share2_reg & x3x4x5x6_second_share ^ x3_share2_reg & x1x4x5x6_second_share ^ x1x3_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x1x3_subscript0_share2_reg ^x4x5_share2_reg & x1x3x6_subscript0_share2_reg ^x4x6_share2_reg & x1x3x5_subscript0_share2_reg ^x5x6_share2_reg & x1x3x4_subscript0_share2_reg ^x6_share2_reg & x1x3x4x5_subscript0_share2_reg ^x5_share2_reg & x1x3x4x6_subscript0_share2_reg ^x4_share2_reg & x1x3x5x6_subscript0_share2_reg ^x1x3x4x5x6_subscript0_share2_reg ;
assign x1x3x4x5x7_second_share =x1_share2_reg & x3x4x5x7_second_share ^ x3_share2_reg & x1x4x5x7_second_share ^ x1x3_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x1x3_subscript0_share2_reg ^x4x5_share2_reg & x1x3x7_subscript0_share2_reg ^x4x7_share2_reg & x1x3x5_subscript0_share2_reg ^x5x7_share2_reg & x1x3x4_subscript0_share2_reg ^x7_share2_reg & x1x3x4x5_subscript0_share2_reg ^x5_share2_reg & x1x3x4x7_subscript0_share2_reg ^x4_share2_reg & x1x3x5x7_subscript0_share2_reg ^x1x3x4x5x7_subscript0_share2_reg ;
assign x1x3x4x6x7_second_share =x1_share2_reg & x3x4x6x7_second_share ^ x3_share2_reg & x1x4x6x7_second_share ^ x1x3_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x1x3_subscript0_share2_reg ^x4x6_share2_reg & x1x3x7_subscript0_share2_reg ^x4x7_share2_reg & x1x3x6_subscript0_share2_reg ^x6x7_share2_reg & x1x3x4_subscript0_share2_reg ^x7_share2_reg & x1x3x4x6_subscript0_share2_reg ^x6_share2_reg & x1x3x4x7_subscript0_share2_reg ^x4_share2_reg & x1x3x6x7_subscript0_share2_reg ^x1x3x4x6x7_subscript0_share2_reg ;
assign x1x3x5x6x7_second_share =x1_share2_reg & x3x5x6x7_second_share ^ x3_share2_reg & x1x5x6x7_second_share ^ x1x3_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x1x3_subscript0_share2_reg ^x5x6_share2_reg & x1x3x7_subscript0_share2_reg ^x5x7_share2_reg & x1x3x6_subscript0_share2_reg ^x6x7_share2_reg & x1x3x5_subscript0_share2_reg ^x7_share2_reg & x1x3x5x6_subscript0_share2_reg ^x6_share2_reg & x1x3x5x7_subscript0_share2_reg ^x5_share2_reg & x1x3x6x7_subscript0_share2_reg ^x1x3x5x6x7_subscript0_share2_reg ;
assign x1x4x5x6x7_second_share =x1_share2_reg & x4x5x6x7_second_share ^ x4_share2_reg & x1x5x6x7_second_share ^ x1x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x1x4_subscript0_share2_reg ^x5x6_share2_reg & x1x4x7_subscript0_share2_reg ^x5x7_share2_reg & x1x4x6_subscript0_share2_reg ^x6x7_share2_reg & x1x4x5_subscript0_share2_reg ^x7_share2_reg & x1x4x5x6_subscript0_share2_reg ^x6_share2_reg & x1x4x5x7_subscript0_share2_reg ^x5_share2_reg & x1x4x6x7_subscript0_share2_reg ^x1x4x5x6x7_subscript0_share2_reg ;
assign x2x3x4x5x6_second_share =x2_share2_reg & x3x4x5x6_second_share ^ x3_share2_reg & x2x4x5x6_second_share ^ x2x3_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x2x3_subscript0_share2_reg ^x4x5_share2_reg & x2x3x6_subscript0_share2_reg ^x4x6_share2_reg & x2x3x5_subscript0_share2_reg ^x5x6_share2_reg & x2x3x4_subscript0_share2_reg ^x6_share2_reg & x2x3x4x5_subscript0_share2_reg ^x5_share2_reg & x2x3x4x6_subscript0_share2_reg ^x4_share2_reg & x2x3x5x6_subscript0_share2_reg ^x2x3x4x5x6_subscript0_share2_reg ;
assign x2x3x4x5x7_second_share =x2_share2_reg & x3x4x5x7_second_share ^ x3_share2_reg & x2x4x5x7_second_share ^ x2x3_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x2x3_subscript0_share2_reg ^x4x5_share2_reg & x2x3x7_subscript0_share2_reg ^x4x7_share2_reg & x2x3x5_subscript0_share2_reg ^x5x7_share2_reg & x2x3x4_subscript0_share2_reg ^x7_share2_reg & x2x3x4x5_subscript0_share2_reg ^x5_share2_reg & x2x3x4x7_subscript0_share2_reg ^x4_share2_reg & x2x3x5x7_subscript0_share2_reg ^x2x3x4x5x7_subscript0_share2_reg ;
assign x2x3x4x6x7_second_share =x2_share2_reg & x3x4x6x7_second_share ^ x3_share2_reg & x2x4x6x7_second_share ^ x2x3_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x2x3_subscript0_share2_reg ^x4x6_share2_reg & x2x3x7_subscript0_share2_reg ^x4x7_share2_reg & x2x3x6_subscript0_share2_reg ^x6x7_share2_reg & x2x3x4_subscript0_share2_reg ^x7_share2_reg & x2x3x4x6_subscript0_share2_reg ^x6_share2_reg & x2x3x4x7_subscript0_share2_reg ^x4_share2_reg & x2x3x6x7_subscript0_share2_reg ^x2x3x4x6x7_subscript0_share2_reg ;
assign x2x3x5x6x7_second_share =x2_share2_reg & x3x5x6x7_second_share ^ x3_share2_reg & x2x5x6x7_second_share ^ x2x3_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x2x3_subscript0_share2_reg ^x5x6_share2_reg & x2x3x7_subscript0_share2_reg ^x5x7_share2_reg & x2x3x6_subscript0_share2_reg ^x6x7_share2_reg & x2x3x5_subscript0_share2_reg ^x7_share2_reg & x2x3x5x6_subscript0_share2_reg ^x6_share2_reg & x2x3x5x7_subscript0_share2_reg ^x5_share2_reg & x2x3x6x7_subscript0_share2_reg ^x2x3x5x6x7_subscript0_share2_reg ;
assign x2x4x5x6x7_second_share =x2_share2_reg & x4x5x6x7_second_share ^ x4_share2_reg & x2x5x6x7_second_share ^ x2x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x2x4_subscript0_share2_reg ^x5x6_share2_reg & x2x4x7_subscript0_share2_reg ^x5x7_share2_reg & x2x4x6_subscript0_share2_reg ^x6x7_share2_reg & x2x4x5_subscript0_share2_reg ^x7_share2_reg & x2x4x5x6_subscript0_share2_reg ^x6_share2_reg & x2x4x5x7_subscript0_share2_reg ^x5_share2_reg & x2x4x6x7_subscript0_share2_reg ^x2x4x5x6x7_subscript0_share2_reg ;
assign x3x4x5x6x7_second_share =x3_share2_reg & x4x5x6x7_second_share ^ x4_share2_reg & x3x5x6x7_second_share ^ x3x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x3x4_subscript0_share2_reg ^x5x6_share2_reg & x3x4x7_subscript0_share2_reg ^x5x7_share2_reg & x3x4x6_subscript0_share2_reg ^x6x7_share2_reg & x3x4x5_subscript0_share2_reg ^x7_share2_reg & x3x4x5x6_subscript0_share2_reg ^x6_share2_reg & x3x4x5x7_subscript0_share2_reg ^x5_share2_reg & x3x4x6x7_subscript0_share2_reg ^x3x4x5x6x7_subscript0_share2_reg ;


// second share of Degree-6 terms

assign x0x1x2x3x4x5_second_share =  x0_share2_reg & x1x2x3x4x5_second_share ^ x1_share2_reg & x0x2x3x4x5_second_share ^ x2_share2_reg & x0x1x3x4x5_second_share ^ x0x1_share2_reg & x2x3x4x5_second_share ^ x0x2_share2_reg & x1x3x4x5_second_share ^ x1x2_share2_reg & x0x3x4x5_second_share ^ x0x1x2_share2_reg & x3x4x5_second_share ^ x3x4x5_share2_reg & x0x1x2_subscript0_share2_reg ^ x3x4_share2_reg & x0x1x2x5_subscript0_share2_reg ^ x4x5_share2_reg & x0x1x2x3_subscript0_share2_reg ^ x3x5_share2_reg & x0x1x2x4_subscript0_share2_reg ^ x3_share2_reg & x0x1x2x4x5_subscript0_share2_reg ^ x4_share2_reg & x0x1x2x3x5_subscript0_share2_reg ^ x5_share2_reg & x0x1x2x3x4_subscript0_share2_reg ^ x0x1x2x3x4x5_subscript0_share2_reg ; 
assign x0x1x2x3x4x6_second_share =  x0_share2_reg & x1x2x3x4x6_second_share ^ x1_share2_reg & x0x2x3x4x6_second_share ^ x2_share2_reg & x0x1x3x4x6_second_share ^ x0x1_share2_reg & x2x3x4x6_second_share ^ x0x2_share2_reg & x1x3x4x6_second_share ^ x1x2_share2_reg & x0x3x4x6_second_share ^ x0x1x2_share2_reg & x3x4x6_second_share ^ x3x4x6_share2_reg & x0x1x2_subscript0_share2_reg ^ x3x4_share2_reg & x0x1x2x6_subscript0_share2_reg ^ x4x6_share2_reg & x0x1x2x3_subscript0_share2_reg ^ x3x6_share2_reg & x0x1x2x4_subscript0_share2_reg ^ x3_share2_reg & x0x1x2x4x6_subscript0_share2_reg ^ x4_share2_reg & x0x1x2x3x6_subscript0_share2_reg ^ x6_share2_reg & x0x1x2x3x4_subscript0_share2_reg ^ x0x1x2x3x4x6_subscript0_share2_reg ;
assign x0x1x2x3x4x7_second_share =  x0_share2_reg & x1x2x3x4x7_second_share ^ x1_share2_reg & x0x2x3x4x7_second_share ^ x2_share2_reg & x0x1x3x4x7_second_share ^ x0x1_share2_reg & x2x3x4x7_second_share ^ x0x2_share2_reg & x1x3x4x7_second_share ^ x1x2_share2_reg & x0x3x4x7_second_share ^ x0x1x2_share2_reg & x3x4x7_second_share ^ x3x4x7_share2_reg & x0x1x2_subscript0_share2_reg ^ x3x4_share2_reg & x0x1x2x7_subscript0_share2_reg ^ x4x7_share2_reg & x0x1x2x3_subscript0_share2_reg ^ x3x7_share2_reg & x0x1x2x4_subscript0_share2_reg ^ x3_share2_reg & x0x1x2x4x7_subscript0_share2_reg ^ x4_share2_reg & x0x1x2x3x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x2x3x4_subscript0_share2_reg ^ x0x1x2x3x4x7_subscript0_share2_reg ;
assign x0x1x2x3x5x6_second_share =  x0_share2_reg & x1x2x3x5x6_second_share ^ x1_share2_reg & x0x2x3x5x6_second_share ^ x2_share2_reg & x0x1x3x5x6_second_share ^ x0x1_share2_reg & x2x3x5x6_second_share ^ x0x2_share2_reg & x1x3x5x6_second_share ^ x1x2_share2_reg & x0x3x5x6_second_share ^ x0x1x2_share2_reg & x3x5x6_second_share ^ x3x5x6_share2_reg & x0x1x2_subscript0_share2_reg ^ x3x5_share2_reg & x0x1x2x6_subscript0_share2_reg ^ x5x6_share2_reg & x0x1x2x3_subscript0_share2_reg ^ x3x6_share2_reg & x0x1x2x5_subscript0_share2_reg ^ x3_share2_reg & x0x1x2x5x6_subscript0_share2_reg ^ x5_share2_reg & x0x1x2x3x6_subscript0_share2_reg ^ x6_share2_reg & x0x1x2x3x5_subscript0_share2_reg ^ x0x1x2x3x5x6_subscript0_share2_reg ;
assign x0x1x2x3x5x7_second_share =  x0_share2_reg & x1x2x3x5x7_second_share ^ x1_share2_reg & x0x2x3x5x7_second_share ^ x2_share2_reg & x0x1x3x5x7_second_share ^ x0x1_share2_reg & x2x3x5x7_second_share ^ x0x2_share2_reg & x1x3x5x7_second_share ^ x1x2_share2_reg & x0x3x5x7_second_share ^ x0x1x2_share2_reg & x3x5x7_second_share ^ x3x5x7_share2_reg & x0x1x2_subscript0_share2_reg ^ x3x5_share2_reg & x0x1x2x7_subscript0_share2_reg ^ x5x7_share2_reg & x0x1x2x3_subscript0_share2_reg ^ x3x7_share2_reg & x0x1x2x5_subscript0_share2_reg ^ x3_share2_reg & x0x1x2x5x7_subscript0_share2_reg ^ x5_share2_reg & x0x1x2x3x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x2x3x5_subscript0_share2_reg ^ x0x1x2x3x5x7_subscript0_share2_reg ;
assign x0x1x2x3x6x7_second_share =  x0_share2_reg & x1x2x3x6x7_second_share ^ x1_share2_reg & x0x2x3x6x7_second_share ^ x2_share2_reg & x0x1x3x6x7_second_share ^ x0x1_share2_reg & x2x3x6x7_second_share ^ x0x2_share2_reg & x1x3x6x7_second_share ^ x1x2_share2_reg & x0x3x6x7_second_share ^ x0x1x2_share2_reg & x3x6x7_second_share ^ x3x6x7_share2_reg & x0x1x2_subscript0_share2_reg ^ x3x6_share2_reg & x0x1x2x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x1x2x3_subscript0_share2_reg ^ x3x7_share2_reg & x0x1x2x6_subscript0_share2_reg ^ x3_share2_reg & x0x1x2x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x1x2x3x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x2x3x6_subscript0_share2_reg ^ x0x1x2x3x6x7_subscript0_share2_reg ;
assign x0x1x2x4x5x6_second_share =  x0_share2_reg & x1x2x4x5x6_second_share ^ x1_share2_reg & x0x2x4x5x6_second_share ^ x2_share2_reg & x0x1x4x5x6_second_share ^ x0x1_share2_reg & x2x4x5x6_second_share ^ x0x2_share2_reg & x1x4x5x6_second_share ^ x1x2_share2_reg & x0x4x5x6_second_share ^ x0x1x2_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x0x1x2_subscript0_share2_reg ^ x4x5_share2_reg & x0x1x2x6_subscript0_share2_reg ^ x5x6_share2_reg & x0x1x2x4_subscript0_share2_reg ^ x4x6_share2_reg & x0x1x2x5_subscript0_share2_reg ^ x4_share2_reg & x0x1x2x5x6_subscript0_share2_reg ^ x5_share2_reg & x0x1x2x4x6_subscript0_share2_reg ^ x6_share2_reg & x0x1x2x4x5_subscript0_share2_reg ^ x0x1x2x4x5x6_subscript0_share2_reg ;
assign x0x1x2x4x5x7_second_share =  x0_share2_reg & x1x2x4x5x7_second_share ^ x1_share2_reg & x0x2x4x5x7_second_share ^ x2_share2_reg & x0x1x4x5x7_second_share ^ x0x1_share2_reg & x2x4x5x7_second_share ^ x0x2_share2_reg & x1x4x5x7_second_share ^ x1x2_share2_reg & x0x4x5x7_second_share ^ x0x1x2_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x0x1x2_subscript0_share2_reg ^ x4x5_share2_reg & x0x1x2x7_subscript0_share2_reg ^ x5x7_share2_reg & x0x1x2x4_subscript0_share2_reg ^ x4x7_share2_reg & x0x1x2x5_subscript0_share2_reg ^ x4_share2_reg & x0x1x2x5x7_subscript0_share2_reg ^ x5_share2_reg & x0x1x2x4x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x2x4x5_subscript0_share2_reg ^ x0x1x2x4x5x7_subscript0_share2_reg ;
assign x0x1x2x4x6x7_second_share =  x0_share2_reg & x1x2x4x6x7_second_share ^ x1_share2_reg & x0x2x4x6x7_second_share ^ x2_share2_reg & x0x1x4x6x7_second_share ^ x0x1_share2_reg & x2x4x6x7_second_share ^ x0x2_share2_reg & x1x4x6x7_second_share ^ x1x2_share2_reg & x0x4x6x7_second_share ^ x0x1x2_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x0x1x2_subscript0_share2_reg ^ x4x6_share2_reg & x0x1x2x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x1x2x4_subscript0_share2_reg ^ x4x7_share2_reg & x0x1x2x6_subscript0_share2_reg ^ x4_share2_reg & x0x1x2x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x1x2x4x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x2x4x6_subscript0_share2_reg ^ x0x1x2x4x6x7_subscript0_share2_reg ;
assign x0x1x2x5x6x7_second_share =  x0_share2_reg & x1x2x5x6x7_second_share ^ x1_share2_reg & x0x2x5x6x7_second_share ^ x2_share2_reg & x0x1x5x6x7_second_share ^ x0x1_share2_reg & x2x5x6x7_second_share ^ x0x2_share2_reg & x1x5x6x7_second_share ^ x1x2_share2_reg & x0x5x6x7_second_share ^ x0x1x2_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x1x2_subscript0_share2_reg ^ x5x6_share2_reg & x0x1x2x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x1x2x5_subscript0_share2_reg ^ x5x7_share2_reg & x0x1x2x6_subscript0_share2_reg ^ x5_share2_reg & x0x1x2x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x1x2x5x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x2x5x6_subscript0_share2_reg ^ x0x1x2x5x6x7_subscript0_share2_reg ;
assign x0x1x3x4x5x6_second_share =  x0_share2_reg & x1x3x4x5x6_second_share ^ x1_share2_reg & x0x3x4x5x6_second_share ^ x3_share2_reg & x0x1x4x5x6_second_share ^ x0x1_share2_reg & x3x4x5x6_second_share ^ x0x3_share2_reg & x1x4x5x6_second_share ^ x1x3_share2_reg & x0x4x5x6_second_share ^ x0x1x3_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x0x1x3_subscript0_share2_reg ^ x4x5_share2_reg & x0x1x3x6_subscript0_share2_reg ^ x5x6_share2_reg & x0x1x3x4_subscript0_share2_reg ^ x4x6_share2_reg & x0x1x3x5_subscript0_share2_reg ^ x4_share2_reg & x0x1x3x5x6_subscript0_share2_reg ^ x5_share2_reg & x0x1x3x4x6_subscript0_share2_reg ^ x6_share2_reg & x0x1x3x4x5_subscript0_share2_reg ^ x0x1x3x4x5x6_subscript0_share2_reg ;
assign x0x1x3x4x5x7_second_share =  x0_share2_reg & x1x3x4x5x7_second_share ^ x1_share2_reg & x0x3x4x5x7_second_share ^ x3_share2_reg & x0x1x4x5x7_second_share ^ x0x1_share2_reg & x3x4x5x7_second_share ^ x0x3_share2_reg & x1x4x5x7_second_share ^ x1x3_share2_reg & x0x4x5x7_second_share ^ x0x1x3_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x0x1x3_subscript0_share2_reg ^ x4x5_share2_reg & x0x1x3x7_subscript0_share2_reg ^ x5x7_share2_reg & x0x1x3x4_subscript0_share2_reg ^ x4x7_share2_reg & x0x1x3x5_subscript0_share2_reg ^ x4_share2_reg & x0x1x3x5x7_subscript0_share2_reg ^ x5_share2_reg & x0x1x3x4x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x3x4x5_subscript0_share2_reg ^ x0x1x3x4x5x7_subscript0_share2_reg ;
assign x0x1x3x4x6x7_second_share =  x0_share2_reg & x1x3x4x6x7_second_share ^ x1_share2_reg & x0x3x4x6x7_second_share ^ x3_share2_reg & x0x1x4x6x7_second_share ^ x0x1_share2_reg & x3x4x6x7_second_share ^ x0x3_share2_reg & x1x4x6x7_second_share ^ x1x3_share2_reg & x0x4x6x7_second_share ^ x0x1x3_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x0x1x3_subscript0_share2_reg ^ x4x6_share2_reg & x0x1x3x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x1x3x4_subscript0_share2_reg ^ x4x7_share2_reg & x0x1x3x6_subscript0_share2_reg ^ x4_share2_reg & x0x1x3x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x1x3x4x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x3x4x6_subscript0_share2_reg ^ x0x1x3x4x6x7_subscript0_share2_reg ;
assign x0x1x3x5x6x7_second_share =  x0_share2_reg & x1x3x5x6x7_second_share ^ x1_share2_reg & x0x3x5x6x7_second_share ^ x3_share2_reg & x0x1x5x6x7_second_share ^ x0x1_share2_reg & x3x5x6x7_second_share ^ x0x3_share2_reg & x1x5x6x7_second_share ^ x1x3_share2_reg & x0x5x6x7_second_share ^ x0x1x3_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x1x3_subscript0_share2_reg ^ x5x6_share2_reg & x0x1x3x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x1x3x5_subscript0_share2_reg ^ x5x7_share2_reg & x0x1x3x6_subscript0_share2_reg ^ x5_share2_reg & x0x1x3x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x1x3x5x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x3x5x6_subscript0_share2_reg ^ x0x1x3x5x6x7_subscript0_share2_reg ;
assign x0x1x4x5x6x7_second_share =  x0_share2_reg & x1x4x5x6x7_second_share ^ x1_share2_reg & x0x4x5x6x7_second_share ^ x4_share2_reg & x0x1x5x6x7_second_share ^ x0x1_share2_reg & x4x5x6x7_second_share ^ x0x4_share2_reg & x1x5x6x7_second_share ^ x1x4_share2_reg & x0x5x6x7_second_share ^ x0x1x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x1x4_subscript0_share2_reg ^ x5x6_share2_reg & x0x1x4x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x1x4x5_subscript0_share2_reg ^ x5x7_share2_reg & x0x1x4x6_subscript0_share2_reg ^ x5_share2_reg & x0x1x4x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x1x4x5x7_subscript0_share2_reg ^ x7_share2_reg & x0x1x4x5x6_subscript0_share2_reg ^ x0x1x4x5x6x7_subscript0_share2_reg ;
assign x0x2x3x4x5x6_second_share =  x0_share2_reg & x2x3x4x5x6_second_share ^ x2_share2_reg & x0x3x4x5x6_second_share ^ x3_share2_reg & x0x2x4x5x6_second_share ^ x0x2_share2_reg & x3x4x5x6_second_share ^ x0x3_share2_reg & x2x4x5x6_second_share ^ x2x3_share2_reg & x0x4x5x6_second_share ^ x0x2x3_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x0x2x3_subscript0_share2_reg ^ x4x5_share2_reg & x0x2x3x6_subscript0_share2_reg ^ x5x6_share2_reg & x0x2x3x4_subscript0_share2_reg ^ x4x6_share2_reg & x0x2x3x5_subscript0_share2_reg ^ x4_share2_reg & x0x2x3x5x6_subscript0_share2_reg ^ x5_share2_reg & x0x2x3x4x6_subscript0_share2_reg ^ x6_share2_reg & x0x2x3x4x5_subscript0_share2_reg ^ x0x2x3x4x5x6_subscript0_share2_reg ;
assign x0x2x3x4x5x7_second_share =  x0_share2_reg & x2x3x4x5x7_second_share ^ x2_share2_reg & x0x3x4x5x7_second_share ^ x3_share2_reg & x0x2x4x5x7_second_share ^ x0x2_share2_reg & x3x4x5x7_second_share ^ x0x3_share2_reg & x2x4x5x7_second_share ^ x2x3_share2_reg & x0x4x5x7_second_share ^ x0x2x3_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x0x2x3_subscript0_share2_reg ^ x4x5_share2_reg & x0x2x3x7_subscript0_share2_reg ^ x5x7_share2_reg & x0x2x3x4_subscript0_share2_reg ^ x4x7_share2_reg & x0x2x3x5_subscript0_share2_reg ^ x4_share2_reg & x0x2x3x5x7_subscript0_share2_reg ^ x5_share2_reg & x0x2x3x4x7_subscript0_share2_reg ^ x7_share2_reg & x0x2x3x4x5_subscript0_share2_reg ^ x0x2x3x4x5x7_subscript0_share2_reg ;
assign x0x2x3x4x6x7_second_share =  x0_share2_reg & x2x3x4x6x7_second_share ^ x2_share2_reg & x0x3x4x6x7_second_share ^ x3_share2_reg & x0x2x4x6x7_second_share ^ x0x2_share2_reg & x3x4x6x7_second_share ^ x0x3_share2_reg & x2x4x6x7_second_share ^ x2x3_share2_reg & x0x4x6x7_second_share ^ x0x2x3_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x0x2x3_subscript0_share2_reg ^ x4x6_share2_reg & x0x2x3x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x2x3x4_subscript0_share2_reg ^ x4x7_share2_reg & x0x2x3x6_subscript0_share2_reg ^ x4_share2_reg & x0x2x3x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x2x3x4x7_subscript0_share2_reg ^ x7_share2_reg & x0x2x3x4x6_subscript0_share2_reg ^ x0x2x3x4x6x7_subscript0_share2_reg ;
assign x0x2x3x5x6x7_second_share =  x0_share2_reg & x2x3x5x6x7_second_share ^ x2_share2_reg & x0x3x5x6x7_second_share ^ x3_share2_reg & x0x2x5x6x7_second_share ^ x0x2_share2_reg & x3x5x6x7_second_share ^ x0x3_share2_reg & x2x5x6x7_second_share ^ x2x3_share2_reg & x0x5x6x7_second_share ^ x0x2x3_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x2x3_subscript0_share2_reg ^ x5x6_share2_reg & x0x2x3x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x2x3x5_subscript0_share2_reg ^ x5x7_share2_reg & x0x2x3x6_subscript0_share2_reg ^ x5_share2_reg & x0x2x3x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x2x3x5x7_subscript0_share2_reg ^ x7_share2_reg & x0x2x3x5x6_subscript0_share2_reg ^ x0x2x3x5x6x7_subscript0_share2_reg ;
assign x0x2x4x5x6x7_second_share =  x0_share2_reg & x2x4x5x6x7_second_share ^ x2_share2_reg & x0x4x5x6x7_second_share ^ x4_share2_reg & x0x2x5x6x7_second_share ^ x0x2_share2_reg & x4x5x6x7_second_share ^ x0x4_share2_reg & x2x5x6x7_second_share ^ x2x4_share2_reg & x0x5x6x7_second_share ^ x0x2x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x2x4_subscript0_share2_reg ^ x5x6_share2_reg & x0x2x4x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x2x4x5_subscript0_share2_reg ^ x5x7_share2_reg & x0x2x4x6_subscript0_share2_reg ^ x5_share2_reg & x0x2x4x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x2x4x5x7_subscript0_share2_reg ^ x7_share2_reg & x0x2x4x5x6_subscript0_share2_reg ^ x0x2x4x5x6x7_subscript0_share2_reg ;
assign x0x3x4x5x6x7_second_share =  x0_share2_reg & x3x4x5x6x7_second_share ^ x3_share2_reg & x0x4x5x6x7_second_share ^ x4_share2_reg & x0x3x5x6x7_second_share ^ x0x3_share2_reg & x4x5x6x7_second_share ^ x0x4_share2_reg & x3x5x6x7_second_share ^ x3x4_share2_reg & x0x5x6x7_second_share ^ x0x3x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x0x3x4_subscript0_share2_reg ^ x5x6_share2_reg & x0x3x4x7_subscript0_share2_reg ^ x6x7_share2_reg & x0x3x4x5_subscript0_share2_reg ^ x5x7_share2_reg & x0x3x4x6_subscript0_share2_reg ^ x5_share2_reg & x0x3x4x6x7_subscript0_share2_reg ^ x6_share2_reg & x0x3x4x5x7_subscript0_share2_reg ^ x7_share2_reg & x0x3x4x5x6_subscript0_share2_reg ^ x0x3x4x5x6x7_subscript0_share2_reg ;
assign x1x2x3x4x5x6_second_share =  x1_share2_reg & x2x3x4x5x6_second_share ^ x2_share2_reg & x1x3x4x5x6_second_share ^ x3_share2_reg & x1x2x4x5x6_second_share ^ x1x2_share2_reg & x3x4x5x6_second_share ^ x1x3_share2_reg & x2x4x5x6_second_share ^ x2x3_share2_reg & x1x4x5x6_second_share ^ x1x2x3_share2_reg & x4x5x6_second_share ^ x4x5x6_share2_reg & x1x2x3_subscript0_share2_reg ^ x4x5_share2_reg & x1x2x3x6_subscript0_share2_reg ^ x5x6_share2_reg & x1x2x3x4_subscript0_share2_reg ^ x4x6_share2_reg & x1x2x3x5_subscript0_share2_reg ^ x4_share2_reg & x1x2x3x5x6_subscript0_share2_reg ^ x5_share2_reg & x1x2x3x4x6_subscript0_share2_reg ^ x6_share2_reg & x1x2x3x4x5_subscript0_share2_reg ^ x1x2x3x4x5x6_subscript0_share2_reg ;
assign x1x2x3x4x5x7_second_share =  x1_share2_reg & x2x3x4x5x7_second_share ^ x2_share2_reg & x1x3x4x5x7_second_share ^ x3_share2_reg & x1x2x4x5x7_second_share ^ x1x2_share2_reg & x3x4x5x7_second_share ^ x1x3_share2_reg & x2x4x5x7_second_share ^ x2x3_share2_reg & x1x4x5x7_second_share ^ x1x2x3_share2_reg & x4x5x7_second_share ^ x4x5x7_share2_reg & x1x2x3_subscript0_share2_reg ^ x4x5_share2_reg & x1x2x3x7_subscript0_share2_reg ^ x5x7_share2_reg & x1x2x3x4_subscript0_share2_reg ^ x4x7_share2_reg & x1x2x3x5_subscript0_share2_reg ^ x4_share2_reg & x1x2x3x5x7_subscript0_share2_reg ^ x5_share2_reg & x1x2x3x4x7_subscript0_share2_reg ^ x7_share2_reg & x1x2x3x4x5_subscript0_share2_reg ^ x1x2x3x4x5x7_subscript0_share2_reg ;
assign x1x2x3x4x6x7_second_share =  x1_share2_reg & x2x3x4x6x7_second_share ^ x2_share2_reg & x1x3x4x6x7_second_share ^ x3_share2_reg & x1x2x4x6x7_second_share ^ x1x2_share2_reg & x3x4x6x7_second_share ^ x1x3_share2_reg & x2x4x6x7_second_share ^ x2x3_share2_reg & x1x4x6x7_second_share ^ x1x2x3_share2_reg & x4x6x7_second_share ^ x4x6x7_share2_reg & x1x2x3_subscript0_share2_reg ^ x4x6_share2_reg & x1x2x3x7_subscript0_share2_reg ^ x6x7_share2_reg & x1x2x3x4_subscript0_share2_reg ^ x4x7_share2_reg & x1x2x3x6_subscript0_share2_reg ^ x4_share2_reg & x1x2x3x6x7_subscript0_share2_reg ^ x6_share2_reg & x1x2x3x4x7_subscript0_share2_reg ^ x7_share2_reg & x1x2x3x4x6_subscript0_share2_reg ^ x1x2x3x4x6x7_subscript0_share2_reg ;
assign x1x2x3x5x6x7_second_share =  x1_share2_reg & x2x3x5x6x7_second_share ^ x2_share2_reg & x1x3x5x6x7_second_share ^ x3_share2_reg & x1x2x5x6x7_second_share ^ x1x2_share2_reg & x3x5x6x7_second_share ^ x1x3_share2_reg & x2x5x6x7_second_share ^ x2x3_share2_reg & x1x5x6x7_second_share ^ x1x2x3_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x1x2x3_subscript0_share2_reg ^ x5x6_share2_reg & x1x2x3x7_subscript0_share2_reg ^ x6x7_share2_reg & x1x2x3x5_subscript0_share2_reg ^ x5x7_share2_reg & x1x2x3x6_subscript0_share2_reg ^ x5_share2_reg & x1x2x3x6x7_subscript0_share2_reg ^ x6_share2_reg & x1x2x3x5x7_subscript0_share2_reg ^ x7_share2_reg & x1x2x3x5x6_subscript0_share2_reg ^ x1x2x3x5x6x7_subscript0_share2_reg ;
assign x1x2x4x5x6x7_second_share =  x1_share2_reg & x2x4x5x6x7_second_share ^ x2_share2_reg & x1x4x5x6x7_second_share ^ x4_share2_reg & x1x2x5x6x7_second_share ^ x1x2_share2_reg & x4x5x6x7_second_share ^ x1x4_share2_reg & x2x5x6x7_second_share ^ x2x4_share2_reg & x1x5x6x7_second_share ^ x1x2x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x1x2x4_subscript0_share2_reg ^ x5x6_share2_reg & x1x2x4x7_subscript0_share2_reg ^ x6x7_share2_reg & x1x2x4x5_subscript0_share2_reg ^ x5x7_share2_reg & x1x2x4x6_subscript0_share2_reg ^ x5_share2_reg & x1x2x4x6x7_subscript0_share2_reg ^ x6_share2_reg & x1x2x4x5x7_subscript0_share2_reg ^ x7_share2_reg & x1x2x4x5x6_subscript0_share2_reg ^ x1x2x4x5x6x7_subscript0_share2_reg ;
assign x1x3x4x5x6x7_second_share =  x1_share2_reg & x3x4x5x6x7_second_share ^ x3_share2_reg & x1x4x5x6x7_second_share ^ x4_share2_reg & x1x3x5x6x7_second_share ^ x1x3_share2_reg & x4x5x6x7_second_share ^ x1x4_share2_reg & x3x5x6x7_second_share ^ x3x4_share2_reg & x1x5x6x7_second_share ^ x1x3x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x1x3x4_subscript0_share2_reg ^ x5x6_share2_reg & x1x3x4x7_subscript0_share2_reg ^ x6x7_share2_reg & x1x3x4x5_subscript0_share2_reg ^ x5x7_share2_reg & x1x3x4x6_subscript0_share2_reg ^ x5_share2_reg & x1x3x4x6x7_subscript0_share2_reg ^ x6_share2_reg & x1x3x4x5x7_subscript0_share2_reg ^ x7_share2_reg & x1x3x4x5x6_subscript0_share2_reg ^ x1x3x4x5x6x7_subscript0_share2_reg ;
assign x2x3x4x5x6x7_second_share =  x2_share2_reg & x3x4x5x6x7_second_share ^ x3_share2_reg & x2x4x5x6x7_second_share ^ x4_share2_reg & x2x3x5x6x7_second_share ^ x2x3_share2_reg & x4x5x6x7_second_share ^ x2x4_share2_reg & x3x5x6x7_second_share ^ x3x4_share2_reg & x2x5x6x7_second_share ^ x2x3x4_share2_reg & x5x6x7_second_share ^ x5x6x7_share2_reg & x2x3x4_subscript0_share2_reg ^ x5x6_share2_reg & x2x3x4x7_subscript0_share2_reg ^ x6x7_share2_reg & x2x3x4x5_subscript0_share2_reg ^ x5x7_share2_reg & x2x3x4x6_subscript0_share2_reg ^ x5_share2_reg & x2x3x4x6x7_subscript0_share2_reg ^ x6_share2_reg & x2x3x4x5x7_subscript0_share2_reg ^ x7_share2_reg & x2x3x4x5x6_subscript0_share2_reg ^ x2x3x4x5x6x7_subscript0_share2_reg ;

// second share of Degree-7 terms

assign x0x1x2x3x4x5x6_second_share = x0_share2_reg & x1x2x3x4x5x6_second_share ^ x1_share2_reg & x0x2x3x4x5x6_second_share ^ x2_share2_reg & x0x1x3x4x5x6_second_share ^ x0x1_share2_reg & x2x3x4x5x6_second_share ^ x0x2_share2_reg & x1x3x4x5x6_second_share ^ x1x2_share2_reg & x0x3x4x5x6_second_share ^ x0x1x2_share2_reg & x3x4x5x6_second_share ^ x3x4x5x6_share2_reg & x0x1x2_subscript0_share2_reg ^x3x4x5_share2_reg & x0x1x2x6_subscript0_share2_reg ^x3x4x6_share2_reg & x0x1x2x5_subscript0_share2_reg ^x3x5x6_share2_reg & x0x1x2x4_subscript0_share2_reg ^x4x5x6_share2_reg & x0x1x2x3_subscript0_share2_reg ^x3x4_share2_reg & x0x1x2x5x6_subscript0_share2_reg ^x3x5_share2_reg & x0x1x2x4x6_subscript0_share2_reg ^x3x6_share2_reg & x0x1x2x4x5_subscript0_share2_reg ^x4x5_share2_reg & x0x1x2x3x6_subscript0_share2_reg ^x4x6_share2_reg & x0x1x2x3x5_subscript0_share2_reg ^x5x6_share2_reg & x0x1x2x3x4_subscript0_share2_reg ^x3_share2_reg & x0x1x2x4x5x6_subscript0_share2_reg ^x4_share2_reg & x0x1x2x3x5x6_subscript0_share2_reg ^x5_share2_reg & x0x1x2x3x4x6_subscript0_share2_reg ^x6_share2_reg & x0x1x2x3x4x5_subscript0_share2_reg ^x0x1x2x3x4x5x6_subscript0_share2_reg ;
assign x0x1x2x3x4x5x7_second_share = x0_share2_reg & x1x2x3x4x5x7_second_share ^ x1_share2_reg & x0x2x3x4x5x7_second_share ^ x2_share2_reg & x0x1x3x4x5x7_second_share ^ x0x1_share2_reg & x2x3x4x5x7_second_share ^ x0x2_share2_reg & x1x3x4x5x7_second_share ^ x1x2_share2_reg & x0x3x4x5x7_second_share ^ x0x1x2_share2_reg & x3x4x5x7_second_share ^ x3x4x5x7_share2_reg & x0x1x2_subscript0_share2_reg ^x3x4x5_share2_reg & x0x1x2x7_subscript0_share2_reg ^x3x4x7_share2_reg & x0x1x2x5_subscript0_share2_reg ^x3x5x7_share2_reg & x0x1x2x4_subscript0_share2_reg ^x4x5x7_share2_reg & x0x1x2x3_subscript0_share2_reg ^x3x4_share2_reg & x0x1x2x5x7_subscript0_share2_reg ^x3x5_share2_reg & x0x1x2x4x7_subscript0_share2_reg ^x3x7_share2_reg & x0x1x2x4x5_subscript0_share2_reg ^x4x5_share2_reg & x0x1x2x3x7_subscript0_share2_reg ^x4x7_share2_reg & x0x1x2x3x5_subscript0_share2_reg ^x5x7_share2_reg & x0x1x2x3x4_subscript0_share2_reg ^x3_share2_reg & x0x1x2x4x5x7_subscript0_share2_reg ^x4_share2_reg & x0x1x2x3x5x7_subscript0_share2_reg ^x5_share2_reg & x0x1x2x3x4x7_subscript0_share2_reg ^x7_share2_reg & x0x1x2x3x4x5_subscript0_share2_reg ^x0x1x2x3x4x5x7_subscript0_share2_reg ;
assign x0x1x2x3x4x6x7_second_share = x0_share2_reg & x1x2x3x4x6x7_second_share ^ x1_share2_reg & x0x2x3x4x6x7_second_share ^ x2_share2_reg & x0x1x3x4x6x7_second_share ^ x0x1_share2_reg & x2x3x4x6x7_second_share ^ x0x2_share2_reg & x1x3x4x6x7_second_share ^ x1x2_share2_reg & x0x3x4x6x7_second_share ^ x0x1x2_share2_reg & x3x4x6x7_second_share ^ x3x4x6x7_share2_reg & x0x1x2_subscript0_share2_reg ^x3x4x6_share2_reg & x0x1x2x7_subscript0_share2_reg ^x3x4x7_share2_reg & x0x1x2x6_subscript0_share2_reg ^x3x6x7_share2_reg & x0x1x2x4_subscript0_share2_reg ^x4x6x7_share2_reg & x0x1x2x3_subscript0_share2_reg ^x3x4_share2_reg & x0x1x2x6x7_subscript0_share2_reg ^x3x6_share2_reg & x0x1x2x4x7_subscript0_share2_reg ^x3x7_share2_reg & x0x1x2x4x6_subscript0_share2_reg ^x4x6_share2_reg & x0x1x2x3x7_subscript0_share2_reg ^x4x7_share2_reg & x0x1x2x3x6_subscript0_share2_reg ^x6x7_share2_reg & x0x1x2x3x4_subscript0_share2_reg ^x3_share2_reg & x0x1x2x4x6x7_subscript0_share2_reg ^x4_share2_reg & x0x1x2x3x6x7_subscript0_share2_reg ^x6_share2_reg & x0x1x2x3x4x7_subscript0_share2_reg ^x7_share2_reg & x0x1x2x3x4x6_subscript0_share2_reg ^x0x1x2x3x4x6x7_subscript0_share2_reg ;
assign x0x1x2x3x5x6x7_second_share = x0_share2_reg & x1x2x3x5x6x7_second_share ^ x1_share2_reg & x0x2x3x5x6x7_second_share ^ x2_share2_reg & x0x1x3x5x6x7_second_share ^ x0x1_share2_reg & x2x3x5x6x7_second_share ^ x0x2_share2_reg & x1x3x5x6x7_second_share ^ x1x2_share2_reg & x0x3x5x6x7_second_share ^ x0x1x2_share2_reg & x3x5x6x7_second_share ^ x3x5x6x7_share2_reg & x0x1x2_subscript0_share2_reg ^x3x5x6_share2_reg & x0x1x2x7_subscript0_share2_reg ^x3x5x7_share2_reg & x0x1x2x6_subscript0_share2_reg ^x3x6x7_share2_reg & x0x1x2x5_subscript0_share2_reg ^x5x6x7_share2_reg & x0x1x2x3_subscript0_share2_reg ^x3x5_share2_reg & x0x1x2x6x7_subscript0_share2_reg ^x3x6_share2_reg & x0x1x2x5x7_subscript0_share2_reg ^x3x7_share2_reg & x0x1x2x5x6_subscript0_share2_reg ^x5x6_share2_reg & x0x1x2x3x7_subscript0_share2_reg ^x5x7_share2_reg & x0x1x2x3x6_subscript0_share2_reg ^x6x7_share2_reg & x0x1x2x3x5_subscript0_share2_reg ^x3_share2_reg & x0x1x2x5x6x7_subscript0_share2_reg ^x5_share2_reg & x0x1x2x3x6x7_subscript0_share2_reg ^x6_share2_reg & x0x1x2x3x5x7_subscript0_share2_reg ^x7_share2_reg & x0x1x2x3x5x6_subscript0_share2_reg ^x0x1x2x3x5x6x7_subscript0_share2_reg ;
assign x0x1x2x4x5x6x7_second_share = x0_share2_reg & x1x2x4x5x6x7_second_share ^ x1_share2_reg & x0x2x4x5x6x7_second_share ^ x2_share2_reg & x0x1x4x5x6x7_second_share ^ x0x1_share2_reg & x2x4x5x6x7_second_share ^ x0x2_share2_reg & x1x4x5x6x7_second_share ^ x1x2_share2_reg & x0x4x5x6x7_second_share ^ x0x1x2_share2_reg & x4x5x6x7_second_share ^ x4x5x6x7_share2_reg & x0x1x2_subscript0_share2_reg ^x4x5x6_share2_reg & x0x1x2x7_subscript0_share2_reg ^x4x5x7_share2_reg & x0x1x2x6_subscript0_share2_reg ^x4x6x7_share2_reg & x0x1x2x5_subscript0_share2_reg ^x5x6x7_share2_reg & x0x1x2x4_subscript0_share2_reg ^x4x5_share2_reg & x0x1x2x6x7_subscript0_share2_reg ^x4x6_share2_reg & x0x1x2x5x7_subscript0_share2_reg ^x4x7_share2_reg & x0x1x2x5x6_subscript0_share2_reg ^x5x6_share2_reg & x0x1x2x4x7_subscript0_share2_reg ^x5x7_share2_reg & x0x1x2x4x6_subscript0_share2_reg ^x6x7_share2_reg & x0x1x2x4x5_subscript0_share2_reg ^x4_share2_reg & x0x1x2x5x6x7_subscript0_share2_reg ^x5_share2_reg & x0x1x2x4x6x7_subscript0_share2_reg ^x6_share2_reg & x0x1x2x4x5x7_subscript0_share2_reg ^x7_share2_reg & x0x1x2x4x5x6_subscript0_share2_reg ^x0x1x2x4x5x6x7_subscript0_share2_reg ;
assign x0x1x3x4x5x6x7_second_share = x0_share2_reg & x1x3x4x5x6x7_second_share ^ x1_share2_reg & x0x3x4x5x6x7_second_share ^ x3_share2_reg & x0x1x4x5x6x7_second_share ^ x0x1_share2_reg & x3x4x5x6x7_second_share ^ x0x3_share2_reg & x1x4x5x6x7_second_share ^ x1x3_share2_reg & x0x4x5x6x7_second_share ^ x0x1x3_share2_reg & x4x5x6x7_second_share ^ x4x5x6x7_share2_reg & x0x1x3_subscript0_share2_reg ^x4x5x6_share2_reg & x0x1x3x7_subscript0_share2_reg ^x4x5x7_share2_reg & x0x1x3x6_subscript0_share2_reg ^x4x6x7_share2_reg & x0x1x3x5_subscript0_share2_reg ^x5x6x7_share2_reg & x0x1x3x4_subscript0_share2_reg ^x4x5_share2_reg & x0x1x3x6x7_subscript0_share2_reg ^x4x6_share2_reg & x0x1x3x5x7_subscript0_share2_reg ^x4x7_share2_reg & x0x1x3x5x6_subscript0_share2_reg ^x5x6_share2_reg & x0x1x3x4x7_subscript0_share2_reg ^x5x7_share2_reg & x0x1x3x4x6_subscript0_share2_reg ^x6x7_share2_reg & x0x1x3x4x5_subscript0_share2_reg ^x4_share2_reg & x0x1x3x5x6x7_subscript0_share2_reg ^x5_share2_reg & x0x1x3x4x6x7_subscript0_share2_reg ^x6_share2_reg & x0x1x3x4x5x7_subscript0_share2_reg ^x7_share2_reg & x0x1x3x4x5x6_subscript0_share2_reg ^x0x1x3x4x5x6x7_subscript0_share2_reg ;
assign x0x2x3x4x5x6x7_second_share = x0_share2_reg & x2x3x4x5x6x7_second_share ^ x2_share2_reg & x0x3x4x5x6x7_second_share ^ x3_share2_reg & x0x2x4x5x6x7_second_share ^ x0x2_share2_reg & x3x4x5x6x7_second_share ^ x0x3_share2_reg & x2x4x5x6x7_second_share ^ x2x3_share2_reg & x0x4x5x6x7_second_share ^ x0x2x3_share2_reg & x4x5x6x7_second_share ^ x4x5x6x7_share2_reg & x0x2x3_subscript0_share2_reg ^x4x5x6_share2_reg & x0x2x3x7_subscript0_share2_reg ^x4x5x7_share2_reg & x0x2x3x6_subscript0_share2_reg ^x4x6x7_share2_reg & x0x2x3x5_subscript0_share2_reg ^x5x6x7_share2_reg & x0x2x3x4_subscript0_share2_reg ^x4x5_share2_reg & x0x2x3x6x7_subscript0_share2_reg ^x4x6_share2_reg & x0x2x3x5x7_subscript0_share2_reg ^x4x7_share2_reg & x0x2x3x5x6_subscript0_share2_reg ^x5x6_share2_reg & x0x2x3x4x7_subscript0_share2_reg ^x5x7_share2_reg & x0x2x3x4x6_subscript0_share2_reg ^x6x7_share2_reg & x0x2x3x4x5_subscript0_share2_reg ^x4_share2_reg & x0x2x3x5x6x7_subscript0_share2_reg ^x5_share2_reg & x0x2x3x4x6x7_subscript0_share2_reg ^x6_share2_reg & x0x2x3x4x5x7_subscript0_share2_reg ^x7_share2_reg & x0x2x3x4x5x6_subscript0_share2_reg ^x0x2x3x4x5x6x7_subscript0_share2_reg ;
assign x1x2x3x4x5x6x7_second_share = x1_share2_reg & x2x3x4x5x6x7_second_share ^ x2_share2_reg & x1x3x4x5x6x7_second_share ^ x3_share2_reg & x1x2x4x5x6x7_second_share ^ x1x2_share2_reg & x3x4x5x6x7_second_share ^ x1x3_share2_reg & x2x4x5x6x7_second_share ^ x2x3_share2_reg & x1x4x5x6x7_second_share ^ x1x2x3_share2_reg & x4x5x6x7_second_share ^ x4x5x6x7_share2_reg & x1x2x3_subscript0_share2_reg ^x4x5x6_share2_reg & x1x2x3x7_subscript0_share2_reg ^x4x5x7_share2_reg & x1x2x3x6_subscript0_share2_reg ^x4x6x7_share2_reg & x1x2x3x5_subscript0_share2_reg ^x5x6x7_share2_reg & x1x2x3x4_subscript0_share2_reg ^x4x5_share2_reg & x1x2x3x6x7_subscript0_share2_reg ^x4x6_share2_reg & x1x2x3x5x7_subscript0_share2_reg ^x4x7_share2_reg & x1x2x3x5x6_subscript0_share2_reg ^x5x6_share2_reg & x1x2x3x4x7_subscript0_share2_reg ^x5x7_share2_reg & x1x2x3x4x6_subscript0_share2_reg ^x6x7_share2_reg & x1x2x3x4x5_subscript0_share2_reg ^x4_share2_reg & x1x2x3x5x6x7_subscript0_share2_reg ^x5_share2_reg & x1x2x3x4x6x7_subscript0_share2_reg ^x6_share2_reg & x1x2x3x4x5x7_subscript0_share2_reg ^x7_share2_reg & x1x2x3x4x5x6_subscript0_share2_reg ^x1x2x3x4x5x6x7_subscript0_share2_reg ;


assign sbox_out1_share2 =  x0x1x2x3x4x6x7_second_share ^ x0x1x2x3x4x6_second_share ^ x0x1x2x3x4x7_second_share ^ x0x1x2x3x4_second_share ^ x0x1x2x3x5x7_second_share ^ x0x1x2x3x6x7_second_share ^ x0x1x2x3x6_second_share ^ x0x1x2x3x7_second_share ^ x0x1x2x3_second_share ^ x0x1x2x4x5x6x7_second_share ^ x0x1x2x4x5x7_second_share ^ x0x1x2x4x5_second_share ^ x0x1x2x4x7_second_share ^ x0x1x2x5x6x7_second_share ^ x0x1x2x5x7_second_share ^ x0x1x2x5_second_share ^ x0x1x2x6x7_second_share ^ x0x1x2x6_second_share ^ x0x1x2x7_second_share ^ x0x1x3x4x6x7_second_share ^ x0x1x3x4x6_second_share ^ x0x1x3x5x6_second_share ^ x0x1x3x5x7_second_share ^ x0x1x3x6x7_second_share ^ x0x1x4x5x6x7_second_share ^ x0x1x4x5x6_second_share ^ x0x1x4x5_second_share ^ x0x1x4x7_second_share ^ x0x1x4_second_share ^ x0x1x5x6x7_second_share ^ x0x1x6_second_share ^ x0x1x7_second_share ^ x0x1_second_share ^ x0x2x3x4x5x6x7_second_share ^ x0x2x3x4x5x6_second_share ^ x0x2x3x4x5x7_second_share ^ x0x2x3x4x5_second_share ^ x0x2x3x4x6_second_share ^ x0x2x3x5x6x7_second_share ^ x0x2x3x5_second_share ^ x0x2x3x7_second_share ^ x0x2x4x5x7_second_share ^ x0x2x4x5_second_share ^ x0x2x4x6x7_second_share ^ x0x2x4x7_second_share ^ x0x2x4_second_share ^ x0x2x5x6_second_share ^ x0x2x5x7_second_share ^ x0x2x5_second_share ^ x0x2x6_second_share ^ x0x2x7_second_share ^ x0x3x4x5x6_second_share ^ x0x3x4x5x7_second_share ^ x0x3x4x6x7_second_share ^ x0x3x4x6_second_share ^ x0x3x4_second_share ^ x0x3x5x6x7_second_share ^ x0x3x5x6_second_share ^ x0x3x5_second_share ^ x0x3x6_second_share ^ x0x4x5x6_second_share ^ x0x4x5x7_second_share ^ x0x4x6x7_second_share ^ x0x4x6_second_share ^ x0x4x7_second_share ^ x0x4_second_share ^ x0x5_second_share ^ x0x6_second_share ^ x0_second_share ^ x1x2x3x4x6x7_second_share ^ x1x2x3x5x6_second_share ^ x1x2x3x5x7_second_share ^ x1x2x3x5_second_share ^ x1x2x3x6_second_share ^ x1x2x3x7_second_share ^ x1x2x3_second_share ^ x1x2x4x5x6x7_second_share ^ x1x2x4x5x6_second_share ^ x1x2x4x6x7_second_share ^ x1x2x4x6_second_share ^ x1x2x4x7_second_share ^ x1x2x4_second_share ^ x1x2x5x6x7_second_share ^ x1x2x6x7_second_share ^ x1x2x6_second_share ^ x1x2_second_share ^ x1x3x4x5x6x7_second_share ^ x1x3x4x5x7_second_share ^ x1x3x4x6_second_share ^ x1x3x4_second_share ^ x1x3x6x7_second_share ^ x1x3x7_second_share ^ x1x3_second_share ^ x1x4x5x6_second_share ^ x1x4x5x7_second_share ^ x1x4x6_second_share ^ x1x4_second_share ^ x1x5x6x7_second_share ^ x1x5x6_second_share ^ x1x6_second_share ^ x2x3x4x5x6x7_second_share ^ x2x3x4x5x6_second_share ^ x2x3x4x5x7_second_share ^ x2x3x5x7_second_share ^ x2x3x5_second_share ^ x2x3x6x7_second_share ^ x2x3x7_second_share ^ x2x3_second_share ^ x2x4x5x6x7_second_share ^ x2x4x5x6_second_share ^ x2x4x5x7_second_share ^ x2x4x7_second_share ^ x2x4_second_share ^ x2x5x6_second_share ^ x2x5x7_second_share ^ x2x6x7_second_share ^ x2x6_second_share ^ x2x7_second_share ^ x2_second_share ^ x3x4x7_second_share ^ x3x5x6x7_second_share ^ x3x5x7_second_share ^ x3x6x7_second_share ^ x3_second_share ^ x4x5x6_second_share ^ x4x6_second_share ^ x4_second_share ^ x5x6x7_second_share ^ x5x6_second_share ^ x5x7_second_share ^ x6x7_second_share ^ 1'b0 ;
assign sbox_out2_share2 =  x0x1x2x3x4x6x7_second_share ^ x0x1x2x3x4x6_second_share ^ x0x1x2x3x4x7_second_share ^ x0x1x2x3x4_second_share ^ x0x1x2x3x5x6x7_second_share ^ x0x1x2x3x5x6_second_share ^ x0x1x2x3x6_second_share ^ x0x1x2x3x7_second_share ^ x0x1x2x4x5x6x7_second_share ^ x0x1x2x4x5x7_second_share ^ x0x1x2x4x5_second_share ^ x0x1x2x4x6x7_second_share ^ x0x1x2x4x6_second_share ^ x0x1x2x4x7_second_share ^ x0x1x2x5x6x7_second_share ^ x0x1x2x6x7_second_share ^ x0x1x2x6_second_share ^ x0x1x3x4x5x6x7_second_share ^ x0x1x3x4x5x6_second_share ^ x0x1x3x4x6x7_second_share ^ x0x1x3x4x6_second_share ^ x0x1x3x4x7_second_share ^ x0x1x3x4_second_share ^ x0x1x3x5x6_second_share ^ x0x1x3x5x7_second_share ^ x0x1x3x6x7_second_share ^ x0x1x3x6_second_share ^ x0x1x3_second_share ^ x0x1x4x5x6_second_share ^ x0x1x4x5_second_share ^ x0x1x4x7_second_share ^ x0x1x4_second_share ^ x0x1x5x6x7_second_share ^ x0x1x5x6_second_share ^ x0x1x6_second_share ^ x0x1_second_share ^ x0x2x3x4x5x6_second_share ^ x0x2x3x4x5x7_second_share ^ x0x2x3x4x5_second_share ^ x0x2x3x4x6x7_second_share ^ x0x2x3x4x7_second_share ^ x0x2x3x5x6x7_second_share ^ x0x2x3x5x7_second_share ^ x0x2x3x6x7_second_share ^ x0x2x3x6_second_share ^ x0x2x3_second_share ^ x0x2x4x5x6_second_share ^ x0x2x4x5_second_share ^ x0x2x5x6x7_second_share ^ x0x2x5x6_second_share ^ x0x2x7_second_share ^ x0x2_second_share ^ x0x3x4x5x7_second_share ^ x0x3x4x5_second_share ^ x0x3x4x6_second_share ^ x0x3x4_second_share ^ x0x3x5x6x7_second_share ^ x0x3_second_share ^ x0x4x5x6x7_second_share ^ x0x4x5x6_second_share ^ x0x4x5x7_second_share ^ x0x4x5_second_share ^ x0x4x6x7_second_share ^ x0x4x6_second_share ^ x0x4x7_second_share ^ x0x4_second_share ^ x0x5x7_second_share ^ x0x6x7_second_share ^ x0x7_second_share ^ x0_second_share ^ x1x2x3x4x5x6_second_share ^ x1x2x3x4x6x7_second_share ^ x1x2x3x4x6_second_share ^ x1x2x3x5x6x7_second_share ^ x1x2x3x5x6_second_share ^ x1x2x3x5_second_share ^ x1x2x3_second_share ^ x1x2x4x5x6_second_share ^ x1x2x4x7_second_share ^ x1x2x4_second_share ^ x1x2x5x6_second_share ^ x1x2x5x7_second_share ^ x1x2x6x7_second_share ^ x1x3x4x5x6x7_second_share ^ x1x3x4x5x6_second_share ^ x1x3x4x5x7_second_share ^ x1x3x4x5_second_share ^ x1x3x4x7_second_share ^ x1x3x4_second_share ^ x1x3x5x6_second_share ^ x1x3x5x7_second_share ^ x1x3x5_second_share ^ x1x3x6_second_share ^ x1x3x7_second_share ^ x1x3_second_share ^ x1x4x5x7_second_share ^ x1x4x6x7_second_share ^ x1x4x7_second_share ^ x1x4_second_share ^ x1x5x6_second_share ^ x1x7_second_share ^ x2x3x4x5x7_second_share ^ x2x3x4x5_second_share ^ x2x3x4x6x7_second_share ^ x2x3x4x7_second_share ^ x2x3x4_second_share ^ x2x3x5x7_second_share ^ x2x3x5_second_share ^ x2x3x6_second_share ^ x2x3_second_share ^ x2x4x5x6x7_second_share ^ x2x4x5x7_second_share ^ x2x4x6x7_second_share ^ x2x5x7_second_share ^ x2x6x7_second_share ^ x2x6_second_share ^ x2x7_second_share ^ x3x4x5x6_second_share ^ x3x4x5x7_second_share ^ x3x4x6x7_second_share ^ x3x4x6_second_share ^ x3x4x7_second_share ^ x3x5x6_second_share ^ x3x5x7_second_share ^ x3x6x7_second_share ^ x3x7_second_share ^ x3_second_share ^ x4x5_second_share ^ x4x6_second_share ^ x5x6x7_second_share ^ x6_second_share ^ x7_second_share ^ 1'b0 ;
assign sbox_out3_share2 =  x0x1x2x3x4x5_second_share ^ x0x1x2x3x4x6x7_second_share ^ x0x1x2x3x4x6_second_share ^ x0x1x2x3x4x7_second_share ^ x0x1x2x3x4_second_share ^ x0x1x2x3x5x6x7_second_share ^ x0x1x2x3x5x6_second_share ^ x0x1x2x3x5_second_share ^ x0x1x2x3x6_second_share ^ x0x1x2x3x7_second_share ^ x0x1x2x4x5x6_second_share ^ x0x1x2x4x5x7_second_share ^ x0x1x2x4x5_second_share ^ x0x1x2x4x7_second_share ^ x0x1x2x5x7_second_share ^ x0x1x2x5_second_share ^ x0x1x2x6x7_second_share ^ x0x1x2x7_second_share ^ x0x1x3x4x5x6x7_second_share ^ x0x1x3x4x5x7_second_share ^ x0x1x3x4x6x7_second_share ^ x0x1x3x4x6_second_share ^ x0x1x3x4x7_second_share ^ x0x1x3x4_second_share ^ x0x1x3x5x6x7_second_share ^ x0x1x3x5x7_second_share ^ x0x1x3x5_second_share ^ x0x1x3x6x7_second_share ^ x0x1x3x6_second_share ^ x0x1x3_second_share ^ x0x1x4x5x6x7_second_share ^ x0x1x4x6x7_second_share ^ x0x1x4x6_second_share ^ x0x1x4_second_share ^ x0x1x5x6_second_share ^ x0x1x5_second_share ^ x0x1x6_second_share ^ x0x1x7_second_share ^ x0x2x3x4x5x6x7_second_share ^ x0x2x3x4x5x6_second_share ^ x0x2x3x4x6x7_second_share ^ x0x2x3x4x7_second_share ^ x0x2x3x4_second_share ^ x0x2x3x5x6x7_second_share ^ x0x2x3x5x7_second_share ^ x0x2x3x5_second_share ^ x0x2x3x7_second_share ^ x0x2x3_second_share ^ x0x2x4x5x6x7_second_share ^ x0x2x4x5x6_second_share ^ x0x2x4x6_second_share ^ x0x2x4x7_second_share ^ x0x2x4_second_share ^ x0x2x5x6x7_second_share ^ x0x2x5_second_share ^ x0x2x7_second_share ^ x0x2_second_share ^ x0x3x4x5x7_second_share ^ x0x3x4x6_second_share ^ x0x3x4x7_second_share ^ x0x3x4_second_share ^ x0x3x5x6x7_second_share ^ x0x3x5x6_second_share ^ x0x3x5x7_second_share ^ x0x3x5_second_share ^ x0x3x6_second_share ^ x0x3x7_second_share ^ x0x3_second_share ^ x0x4x5x6x7_second_share ^ x0x4x5_second_share ^ x0x4x6_second_share ^ x0x4x7_second_share ^ x0x4_second_share ^ x0x5x7_second_share ^ x0x5_second_share ^ x0x6x7_second_share ^ x0x6_second_share ^ x0x7_second_share ^ x0_second_share ^ x1x2x3x4x5x6x7_second_share ^ x1x2x3x4x5x7_second_share ^ x1x2x3x4x5_second_share ^ x1x2x3x4x6x7_second_share ^ x1x2x3x4x6_second_share ^ x1x2x3x4_second_share ^ x1x2x3x5_second_share ^ x1x2x3x6x7_second_share ^ x1x2x3x6_second_share ^ x1x2x4x5x6_second_share ^ x1x2x4x5x7_second_share ^ x1x2x4x6x7_second_share ^ x1x2x4x7_second_share ^ x1x2x4_second_share ^ x1x2x5x7_second_share ^ x1x2x5_second_share ^ x1x2x6x7_second_share ^ x1x2x6_second_share ^ x1x2x7_second_share ^ x1x3x4x5x6_second_share ^ x1x3x4x6x7_second_share ^ x1x3x4_second_share ^ x1x3x5x6x7_second_share ^ x1x3x5x7_second_share ^ x1x3x5_second_share ^ x1x3x6x7_second_share ^ x1x3x7_second_share ^ x1x4x5x6x7_second_share ^ x1x4x5x7_second_share ^ x1x4x5_second_share ^ x1x4x7_second_share ^ x1x4_second_share ^ x1x5x6x7_second_share ^ x1x5x6_second_share ^ x1x5x7_second_share ^ x1_second_share ^ x2x3x4x5x6x7_second_share ^ x2x3x4x6x7_second_share ^ x2x3x4x6_second_share ^ x2x3x4x7_second_share ^ x2x3x4_second_share ^ x2x3x5x6x7_second_share ^ x2x3x5x6_second_share ^ x2x3x6_second_share ^ x2x3x7_second_share ^ x2x3_second_share ^ x2x4x5x6_second_share ^ x2x4x5x7_second_share ^ x2x4x5_second_share ^ x2x4x6x7_second_share ^ x2x5x6x7_second_share ^ x2x6x7_second_share ^ x3x4x5x6x7_second_share ^ x3x4x5x6_second_share ^ x3x4x5_second_share ^ x3x4x6_second_share ^ x3x4_second_share ^ x3x5x6x7_second_share ^ x3x5x6_second_share ^ x4x5x6x7_second_share ^ x4x6x7_second_share ^ x4x7_second_share ^ x5x6_second_share ^ x5_second_share ^ x6x7_second_share ^ x7_second_share ;
assign sbox_out4_share2 =  x0x1x2x3x4x5x6_second_share ^ x0x1x2x3x4x6_second_share ^ x0x1x2x3x4x7_second_share ^ x0x1x2x3x4_second_share ^ x0x1x2x3x5x6x7_second_share ^ x0x1x2x3x5x6_second_share ^ x0x1x2x3x5x7_second_share ^ x0x1x2x3x5_second_share ^ x0x1x2x3x6x7_second_share ^ x0x1x2x3x7_second_share ^ x0x1x2x3_second_share ^ x0x1x2x4x5x7_second_share ^ x0x1x2x4x6x7_second_share ^ x0x1x2x4x7_second_share ^ x0x1x2x4_second_share ^ x0x1x2x5x6_second_share ^ x0x1x2x5x7_second_share ^ x0x1x2x5_second_share ^ x0x1x3x4x5x6x7_second_share ^ x0x1x3x4x5x7_second_share ^ x0x1x3x4x5_second_share ^ x0x1x3x4x6_second_share ^ x0x1x3x4x7_second_share ^ x0x1x3x5x6_second_share ^ x0x1x3x6_second_share ^ x0x1x3_second_share ^ x0x1x4x5x7_second_share ^ x0x1x4x6_second_share ^ x0x1x4_second_share ^ x0x1x5x6x7_second_share ^ x0x1x5x6_second_share ^ x0x1x5_second_share ^ x0x1x6x7_second_share ^ x0x1x6_second_share ^ x0x1x7_second_share ^ x0x2x3x4x5x6x7_second_share ^ x0x2x3x4x5_second_share ^ x0x2x3x4x6x7_second_share ^ x0x2x3x5x6x7_second_share ^ x0x2x3x5x6_second_share ^ x0x2x3x5x7_second_share ^ x0x2x3x6x7_second_share ^ x0x2x3x7_second_share ^ x0x2x3_second_share ^ x0x2x4x5x6_second_share ^ x0x2x4x5x7_second_share ^ x0x2x4x6_second_share ^ x0x2x4x7_second_share ^ x0x2x4_second_share ^ x0x2x5x6x7_second_share ^ x0x2x5x6_second_share ^ x0x2x6x7_second_share ^ x0x2x6_second_share ^ x0x2x7_second_share ^ x0x3x4x5x6_second_share ^ x0x3x4x5x7_second_share ^ x0x3x4x6x7_second_share ^ x0x3x4x6_second_share ^ x0x3x4_second_share ^ x0x3x5x6x7_second_share ^ x0x3x6x7_second_share ^ x0x3x6_second_share ^ x0x3x7_second_share ^ x0x3_second_share ^ x0x4x5x6x7_second_share ^ x0x4x5x6_second_share ^ x0x4x5_second_share ^ x0x4x6_second_share ^ x0x5x6x7_second_share ^ x0x7_second_share ^ x0_second_share ^ x1x2x3x4x5x6_second_share ^ x1x2x3x4x5x7_second_share ^ x1x2x3x4x6x7_second_share ^ x1x2x3x5x6x7_second_share ^ x1x2x3x5x6_second_share ^ x1x2x3x5_second_share ^ x1x2x3x6_second_share ^ x1x2x3x7_second_share ^ x1x2x3_second_share ^ x1x2x4x5x6x7_second_share ^ x1x2x4x5x6_second_share ^ x1x2x4x5_second_share ^ x1x2x4x7_second_share ^ x1x2x5x6x7_second_share ^ x1x2x5x7_second_share ^ x1x2x5_second_share ^ x1x2x6x7_second_share ^ x1x2x6_second_share ^ x1x2x7_second_share ^ x1x2_second_share ^ x1x3x4x5_second_share ^ x1x3x4x6x7_second_share ^ x1x3x4x6_second_share ^ x1x3x4x7_second_share ^ x1x3x4_second_share ^ x1x3x5x6x7_second_share ^ x1x3x5x6_second_share ^ x1x4x5x6_second_share ^ x1x4x5x7_second_share ^ x1x4x6x7_second_share ^ x1x5x6x7_second_share ^ x1x5x6_second_share ^ x1x7_second_share ^ x2x3x4x5x6x7_second_share ^ x2x3x4x5x6_second_share ^ x2x3x4x5x7_second_share ^ x2x3x4x5_second_share ^ x2x3x4_second_share ^ x2x3x5_second_share ^ x2x3x7_second_share ^ x2x3_second_share ^ x2x4x5x6x7_second_share ^ x2x4x5x6_second_share ^ x2x4x5x7_second_share ^ x2x4x5_second_share ^ x2x4x6x7_second_share ^ x2x5x7_second_share ^ x3x4x5x6x7_second_share ^ x3x4x5x6_second_share ^ x3x4x6x7_second_share ^ x3x4x7_second_share ^ x3x5x6x7_second_share ^ x3x5x6_second_share ^ x3x5x7_second_share ^ x3x6_second_share ^ x3x7_second_share ^ x4x5x6x7_second_share ^ x4x5_second_share ^ x4_second_share ^ x5x6x7_second_share ^ x5x6_second_share ^ x5x7_second_share ^ x6x7_second_share ^ x6_second_share ^ x7_second_share ;
assign sbox_out5_share2 =  x0x1x2x3x4x5x7_second_share ^ x0x1x2x3x4x5_second_share ^ x0x1x2x3x4x6x7_second_share ^ x0x1x2x3x4x7_second_share ^ x0x1x2x3x4_second_share ^ x0x1x2x3x5x6_second_share ^ x0x1x2x3x6_second_share ^ x0x1x2x3x7_second_share ^ x0x1x2x4x5x6_second_share ^ x0x1x2x4x5_second_share ^ x0x1x2x5x7_second_share ^ x0x1x2x6x7_second_share ^ x0x1x2x6_second_share ^ x0x1x3x4x5x6_second_share ^ x0x1x3x4x6_second_share ^ x0x1x3x5x7_second_share ^ x0x1x3x5_second_share ^ x0x1x3x6x7_second_share ^ x0x1x3x6_second_share ^ x0x1x3x7_second_share ^ x0x1x4x5x6_second_share ^ x0x1x4x5_second_share ^ x0x1x4x6_second_share ^ x0x1x5x6x7_second_share ^ x0x1x5x6_second_share ^ x0x1x5x7_second_share ^ x0x1x6x7_second_share ^ x0x1_second_share ^ x0x2x3x4x5x6x7_second_share ^ x0x2x3x4x5x7_second_share ^ x0x2x3x4x5_second_share ^ x0x2x3x4x6_second_share ^ x0x2x3x4_second_share ^ x0x2x3x5x6_second_share ^ x0x2x3x5x7_second_share ^ x0x2x3_second_share ^ x0x2x4x6x7_second_share ^ x0x2x5x7_second_share ^ x0x2x6_second_share ^ x0x3x4x5x6x7_second_share ^ x0x3x4x5_second_share ^ x0x3x4x6x7_second_share ^ x0x3x4x6_second_share ^ x0x3x4x7_second_share ^ x0x3x4_second_share ^ x0x3x5x6x7_second_share ^ x0x3x5x6_second_share ^ x0x3x5x7_second_share ^ x0x3x5_second_share ^ x0x3x6x7_second_share ^ x0x4x5x6x7_second_share ^ x0x4x5x6_second_share ^ x0x4x5_second_share ^ x0x4x6x7_second_share ^ x0x4x6_second_share ^ x0x4x7_second_share ^ x0x4_second_share ^ x0x5_second_share ^ x0x6x7_second_share ^ x0x6_second_share ^ x0x7_second_share ^ x0_second_share ^ x1x2x3x4x5x6_second_share ^ x1x2x3x4x5x7_second_share ^ x1x2x3x4x6x7_second_share ^ x1x2x3x4x6_second_share ^ x1x2x3x4_second_share ^ x1x2x3x5x6x7_second_share ^ x1x2x3x5x6_second_share ^ x1x2x3x5x7_second_share ^ x1x2x3x5_second_share ^ x1x2x4x5x6_second_share ^ x1x2x4x5x7_second_share ^ x1x2x4x6_second_share ^ x1x2x4_second_share ^ x1x2x5x6x7_second_share ^ x1x2x5x7_second_share ^ x1x2x6x7_second_share ^ x1x3x4x5x6_second_share ^ x1x3x4x5x7_second_share ^ x1x3x4x5_second_share ^ x1x3x4x7_second_share ^ x1x3x5x6x7_second_share ^ x1x3x5_second_share ^ x1x4x5x6x7_second_share ^ x1x4x5_second_share ^ x1x4_second_share ^ x1x5x7_second_share ^ x1x5_second_share ^ x1x6x7_second_share ^ x1x6_second_share ^ x1_second_share ^ x2x3x4x5x6_second_share ^ x2x3x4x5x7_second_share ^ x2x3x4x6x7_second_share ^ x2x3x4x7_second_share ^ x2x3x4_second_share ^ x2x3x5x6_second_share ^ x2x3x5x7_second_share ^ x2x3x5_second_share ^ x2x3x6_second_share ^ x2x3_second_share ^ x2x4x5x6x7_second_share ^ x2x4x5_second_share ^ x2x4x7_second_share ^ x2x5x6_second_share ^ x2x5_second_share ^ x2x6x7_second_share ^ x2_second_share ^ x3x4x5x6x7_second_share ^ x3x4x5x7_second_share ^ x3x4x5_second_share ^ x3x4x6x7_second_share ^ x3x4x6_second_share ^ x3x4x7_second_share ^ x3x4_second_share ^ x3x5x6x7_second_share ^ x3x5x6_second_share ^ x3x5x7_second_share ^ x3x5_second_share ^ x3x6x7_second_share ^ x3x7_second_share ^ x3_second_share ^ x4x5x7_second_share ^ x4x5_second_share ^ x4x6x7_second_share ^ x4x6_second_share ^ x5x6x7_second_share ^ x5x7_second_share ^ x5_second_share ^ x6x7_second_share ;
assign sbox_out6_share2 =  x0x1x2x3x4x5_second_share ^ x0x1x2x3x4_second_share ^ x0x1x2x3x5x6x7_second_share ^ x0x1x2x3x5x6_second_share ^ x0x1x2x3x5x7_second_share ^ x0x1x2x3x5_second_share ^ x0x1x2x3x6_second_share ^ x0x1x2x3x7_second_share ^ x0x1x2x3_second_share ^ x0x1x2x4x5x6x7_second_share ^ x0x1x2x4x5x6_second_share ^ x0x1x2x4x5x7_second_share ^ x0x1x2x4x5_second_share ^ x0x1x2x4x6_second_share ^ x0x1x2x5_second_share ^ x0x1x2x6x7_second_share ^ x0x1x2_second_share ^ x0x1x3x4_second_share ^ x0x1x3x5x7_second_share ^ x0x1x3x7_second_share ^ x0x1x3_second_share ^ x0x1x4x5x6_second_share ^ x0x1x4x5x7_second_share ^ x0x1x4x5_second_share ^ x0x1x4x6x7_second_share ^ x0x1x4x6_second_share ^ x0x1x4x7_second_share ^ x0x1x4_second_share ^ x0x1x5x6x7_second_share ^ x0x1x5x6_second_share ^ x0x1x5x7_second_share ^ x0x1x5_second_share ^ x0x1x6_second_share ^ x0x1x7_second_share ^ x0x2x3x4x6x7_second_share ^ x0x2x3x4x7_second_share ^ x0x2x3x4_second_share ^ x0x2x3x5x7_second_share ^ x0x2x3x5_second_share ^ x0x2x3x6x7_second_share ^ x0x2x4x5x6x7_second_share ^ x0x2x4x5x7_second_share ^ x0x2x4x5_second_share ^ x0x2x4_second_share ^ x0x2x6_second_share ^ x0x3x4x5x6_second_share ^ x0x3x4x5x7_second_share ^ x0x3x4x7_second_share ^ x0x3x5_second_share ^ x0x3_second_share ^ x0x4x5x6x7_second_share ^ x0x4x6x7_second_share ^ x0x4x7_second_share ^ x0x5x6x7_second_share ^ x0x5x6_second_share ^ x1x2x3x4x6x7_second_share ^ x1x2x3x4x6_second_share ^ x1x2x3x4x7_second_share ^ x1x2x3x5x6x7_second_share ^ x1x2x3x5_second_share ^ x1x2x3x6_second_share ^ x1x2x4x5x6x7_second_share ^ x1x2x4x5x6_second_share ^ x1x2x4x5_second_share ^ x1x2x4x7_second_share ^ x1x2x4_second_share ^ x1x2x5_second_share ^ x1x2x6_second_share ^ x1x3x4x5x6_second_share ^ x1x3x4x6x7_second_share ^ x1x3x4x6_second_share ^ x1x3x4x7_second_share ^ x1x3x5x6_second_share ^ x1x3x5x7_second_share ^ x1x3x5_second_share ^ x1x3x6_second_share ^ x1x3x7_second_share ^ x1x4x5x7_second_share ^ x1x4x6_second_share ^ x1x4x7_second_share ^ x1x5x6_second_share ^ x1x5x7_second_share ^ x1x5_second_share ^ x1x6x7_second_share ^ x1x6_second_share ^ x2x3x4x5x6_second_share ^ x2x3x4x5_second_share ^ x2x3x4x6_second_share ^ x2x3x4x7_second_share ^ x2x3x5x6x7_second_share ^ x2x3x5x6_second_share ^ x2x3x6_second_share ^ x2x3x7_second_share ^ x2x4x5x6x7_second_share ^ x2x4x5x7_second_share ^ x2x4x5_second_share ^ x2x4x7_second_share ^ x2x4_second_share ^ x2x5x7_second_share ^ x2x6x7_second_share ^ x3x4x5x6_second_share ^ x3x4x5x7_second_share ^ x3x4x5_second_share ^ x3x4x6x7_second_share ^ x3x4_second_share ^ x3x5x7_second_share ^ x4x5x7_second_share ^ x4x6_second_share ^ x4_second_share ^ x5x6x7_second_share ^ x5x7_second_share ^ x6_second_share ^ x7_second_share ^ 1'b0 ;
assign sbox_out7_share2 =  x0x1x2x3x4x7_second_share ^ x0x1x2x3x5x6_second_share ^ x0x1x2x3x5_second_share ^ x0x1x2x3x6_second_share ^ x0x1x2x3x7_second_share ^ x0x1x2x4x5x6x7_second_share ^ x0x1x2x4x5x6_second_share ^ x0x1x2x4x5x7_second_share ^ x0x1x2x4x6x7_second_share ^ x0x1x2x4_second_share ^ x0x1x2x5x6x7_second_share ^ x0x1x2x5_second_share ^ x0x1x3x4x5x6x7_second_share ^ x0x1x3x4x5x6_second_share ^ x0x1x3x4x5x7_second_share ^ x0x1x3x4x5_second_share ^ x0x1x3x4x6x7_second_share ^ x0x1x3x4_second_share ^ x0x1x3x5x6x7_second_share ^ x0x1x3x6x7_second_share ^ x0x1x3x6_second_share ^ x0x1x3x7_second_share ^ x0x1x3_second_share ^ x0x1x4x5x7_second_share ^ x0x1x4_second_share ^ x0x1x5_second_share ^ x0x1x6x7_second_share ^ x0x2x3x4x5_second_share ^ x0x2x3x5x6_second_share ^ x0x2x3x5_second_share ^ x0x2x3x6_second_share ^ x0x2x3x7_second_share ^ x0x2x4x5x7_second_share ^ x0x2x4x5_second_share ^ x0x2x4x6x7_second_share ^ x0x2x4x6_second_share ^ x0x2x4_second_share ^ x0x2x5x6x7_second_share ^ x0x2x5x7_second_share ^ x0x2x5_second_share ^ x0x2x6_second_share ^ x0x3x4x6x7_second_share ^ x0x3x4x6_second_share ^ x0x3x4x7_second_share ^ x0x3x5_second_share ^ x0x3x6_second_share ^ x0x4x5x6x7_second_share ^ x0x4x5_second_share ^ x0x4x6x7_second_share ^ x0x4x6_second_share ^ x0x4x7_second_share ^ x0x4_second_share ^ x0x5x6_second_share ^ x0x5x7_second_share ^ x0x5_second_share ^ x0x7_second_share ^ x1x2x3x4x5_second_share ^ x1x2x3x4x7_second_share ^ x1x2x3x4_second_share ^ x1x2x3x5x7_second_share ^ x1x2x3x5_second_share ^ x1x2x3x6_second_share ^ x1x2x4x5x6_second_share ^ x1x2x4x5_second_share ^ x1x2x4x7_second_share ^ x1x2x5x6x7_second_share ^ x1x2x5_second_share ^ x1x2x6_second_share ^ x1x2x7_second_share ^ x1x3x4x5x6x7_second_share ^ x1x3x4x5x6_second_share ^ x1x3x4x5x7_second_share ^ x1x3x4x6_second_share ^ x1x3x4x7_second_share ^ x1x3x4_second_share ^ x1x3x5x7_second_share ^ x1x3x6_second_share ^ x1x3_second_share ^ x1x4x5x6x7_second_share ^ x1x4x5x7_second_share ^ x1x4x6x7_second_share ^ x1x4x6_second_share ^ x1x4x7_second_share ^ x1x5x6_second_share ^ x1x6x7_second_share ^ x1x7_second_share ^ x2x3x4x5_second_share ^ x2x3x4x6x7_second_share ^ x2x3x4x6_second_share ^ x2x3x4_second_share ^ x2x3x5x6x7_second_share ^ x2x3x5x6_second_share ^ x2x3x5x7_second_share ^ x2x3x7_second_share ^ x2x3_second_share ^ x2x4x6_second_share ^ x2x4x7_second_share ^ x3x4x5x6x7_second_share ^ x3x4x6_second_share ^ x3x5x7_second_share ^ x3x5_second_share ^ x3x6x7_second_share ^ x3x7_second_share ^ x3_second_share ^ x4x5x6x7_second_share ^ x4x5x6_second_share ^ x4x6_second_share ^ x5x6x7_second_share ^ x5x7_second_share ^ x5_second_share ^ x6_second_share ^ 1'b0 ;
assign sbox_out8_share2 =  x0x1x2x3x4_second_share ^ x0x1x2x3x6x7_second_share ^ x0x1x2x3x6_second_share ^ x0x1x2x3_second_share ^ x0x1x2x4x5x7_second_share ^ x0x1x2x4x6_second_share ^ x0x1x2x4_second_share ^ x0x1x2x5x7_second_share ^ x0x1x2x5_second_share ^ x0x1x2x6x7_second_share ^ x0x1x2x7_second_share ^ x0x1x3x4x5x6x7_second_share ^ x0x1x3x4x5x7_second_share ^ x0x1x3x4x5_second_share ^ x0x1x3x4x6x7_second_share ^ x0x1x3x4x7_second_share ^ x0x1x3x4_second_share ^ x0x1x3x5x6x7_second_share ^ x0x1x3x6_second_share ^ x0x1x4x5x6_second_share ^ x0x1x4x5x7_second_share ^ x0x1x4x7_second_share ^ x0x1x4_second_share ^ x0x1x5x6x7_second_share ^ x0x1x5_second_share ^ x0x1x6_second_share ^ x0x2x3x4x5x6x7_second_share ^ x0x2x3x4x5x6_second_share ^ x0x2x3x4x5x7_second_share ^ x0x2x3x4x5_second_share ^ x0x2x3x4x6x7_second_share ^ x0x2x3x4x6_second_share ^ x0x2x3x4x7_second_share ^ x0x2x3x5x6x7_second_share ^ x0x2x3x5_second_share ^ x0x2x3x6_second_share ^ x0x2x3x7_second_share ^ x0x2x3_second_share ^ x0x2x4x5x6x7_second_share ^ x0x2x4x6_second_share ^ x0x2x4x7_second_share ^ x0x2x5_second_share ^ x0x2x7_second_share ^ x0x2_second_share ^ x0x3x4x5x6_second_share ^ x0x3x4x6x7_second_share ^ x0x3x4x6_second_share ^ x0x3x4x7_second_share ^ x0x3x5x6x7_second_share ^ x0x3x5x6_second_share ^ x0x3x5x7_second_share ^ x0x3x5_second_share ^ x0x3x6x7_second_share ^ x0x3x6_second_share ^ x0x3x7_second_share ^ x0x4x5_second_share ^ x0x4x6x7_second_share ^ x0x5x6_second_share ^ x0x6x7_second_share ^ x0x6_second_share ^ x0x7_second_share ^ x1x2x3x4_second_share ^ x1x2x3x5x6_second_share ^ x1x2x3x5_second_share ^ x1x2x3x7_second_share ^ x1x2x3_second_share ^ x1x2x4x5x6_second_share ^ x1x2x4x5_second_share ^ x1x2x4x6x7_second_share ^ x1x2x4x6_second_share ^ x1x2x5x6x7_second_share ^ x1x2x6_second_share ^ x1x2_second_share ^ x1x3x4x5x6x7_second_share ^ x1x3x4x7_second_share ^ x1x3x5x6x7_second_share ^ x1x3x5_second_share ^ x1x3x6x7_second_share ^ x1x3x6_second_share ^ x1x4x5x6x7_second_share ^ x1x4x5x7_second_share ^ x1x4x6x7_second_share ^ x1x4x7_second_share ^ x1x5x6x7_second_share ^ x1x7_second_share ^ x2x3x4x5x6_second_share ^ x2x3x4x7_second_share ^ x2x3x5_second_share ^ x2x4x6x7_second_share ^ x2x4x6_second_share ^ x2x4_second_share ^ x2x5x6x7_second_share ^ x2x5x6_second_share ^ x2x6x7_second_share ^ x2x6_second_share ^ x2_second_share ^ x3x4x5x6x7_second_share ^ x3x4x5x6_second_share ^ x3x4x5_second_share ^ x3x5x7_second_share ^ x3x5_second_share ^ x4x5x6x7_second_share ^ x4x5x6_second_share ^ x4x5x7_second_share ^ x4x6x7_second_share ^ x4x6_second_share ^ x4_second_share ^ x5x7_second_share ^ x5_second_share ^ x7_second_share ;


endmodule